module wisard_lut
#(parameter ADDR_WIDTH=16, INDEX_WIDTH=9, O_WIDTH=10)
(input [ADDR_WIDTH-1:0] addr, input [INDEX_WIDTH-1:0] index, output [O_WIDTH-1:0] out);


reg [9:0] out_v [0:391];


assign out = out_v[index];

always @(*) begin
  case (addr)
    16'b0000010000000000: out_v[0] = 10'b0011101001;
    16'b0000011001010000: out_v[0] = 10'b0110001101;
    16'b0000001001010000: out_v[0] = 10'b0100000101;
    16'b0000001001000000: out_v[0] = 10'b0100010111;
    16'b0000000001000000: out_v[0] = 10'b0100011101;
    16'b0000001000010000: out_v[0] = 10'b0010001001;
    16'b0000001000000000: out_v[0] = 10'b0101011100;
    16'b0000011001000000: out_v[0] = 10'b0010011001;
    16'b0000010001000000: out_v[0] = 10'b1010011011;
    16'b0000000001010000: out_v[0] = 10'b0000010111;
    16'b0000010001010000: out_v[0] = 10'b0111000000;
    16'b0001001001000000: out_v[0] = 10'b0001001010;
    16'b0000001001000100: out_v[0] = 10'b1011110011;
    16'b0000001001110000: out_v[0] = 10'b0110110011;
    16'b0000000001110000: out_v[0] = 10'b0110010001;
    16'b0000000000010000: out_v[0] = 10'b1011011000;
    16'b0001000001000000: out_v[0] = 10'b0100100111;
    16'b0000011000010000: out_v[0] = 10'b0111000000;
    16'b0000001000110000: out_v[0] = 10'b1001100001;
    16'b0000000000000000: out_v[0] = 10'b0110110111;
    16'b0000000001100000: out_v[0] = 10'b0001010000;
    16'b0000000000110000: out_v[0] = 10'b0010111010;
    16'b0001000000000000: out_v[0] = 10'b0001000111;
    16'b0000000000000010: out_v[0] = 10'b1111001101;
    16'b0001000001000010: out_v[0] = 10'b0010000101;
    16'b0001001000000000: out_v[0] = 10'b0010110010;
    16'b0000001101000000: out_v[0] = 10'b0001100111;
    16'b0000000101000000: out_v[0] = 10'b0101011111;
    16'b0000001001000010: out_v[0] = 10'b0111111110;
    16'b0001001101000000: out_v[0] = 10'b1101101011;
    16'b0001001001000010: out_v[0] = 10'b1011111001;
    16'b0000001100000000: out_v[0] = 10'b0011000000;
    16'b0000000001000010: out_v[0] = 10'b1000110110;
    16'b0000010000010000: out_v[0] = 10'b0000101000;
    16'b0000011000000000: out_v[0] = 10'b1010000000;
    16'b1000010000000000: out_v[0] = 10'b0110101000;
    16'b0000011010000000: out_v[0] = 10'b0010110011;
    16'b1000000000000000: out_v[0] = 10'b1111011001;
    16'b0000000010000000: out_v[0] = 10'b1101010000;
    16'b0000000000100000: out_v[0] = 10'b0010101110;
    16'b1000000010000000: out_v[0] = 10'b1010100001;
    16'b0000001001100000: out_v[0] = 10'b1001010010;
    16'b0000001000000100: out_v[0] = 10'b1010011011;
    16'b0000000011000000: out_v[0] = 10'b1001101110;
    16'b0000000000000100: out_v[0] = 10'b1110001010;
    16'b0000001000100000: out_v[0] = 10'b1101110110;
    16'b0000001000000010: out_v[0] = 10'b0101000101;
    16'b1000000000000100: out_v[0] = 10'b1111111111;
    16'b1000001000000000: out_v[0] = 10'b1010000010;
    16'b0000010000000100: out_v[0] = 10'b1001000111;
    16'b1000000010000100: out_v[0] = 10'b0111011010;
    16'b1000000001000000: out_v[0] = 10'b1010100010;
    16'b1000100000000000: out_v[0] = 10'b1101011111;
    16'b0000100000000000: out_v[0] = 10'b1101001110;
    16'b0000110000000000: out_v[0] = 10'b1010110101;
    16'b1000000011000000: out_v[0] = 10'b1001100001;
    default: out_v[0] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000010010110: out_v[1] = 10'b0001001111;
    16'b1000000010010110: out_v[1] = 10'b0110011111;
    16'b1000000010010111: out_v[1] = 10'b1110111110;
    16'b1000000000010111: out_v[1] = 10'b1010011110;
    16'b0000001010010110: out_v[1] = 10'b0001000011;
    16'b1100000000010101: out_v[1] = 10'b0110000001;
    16'b1000000010010101: out_v[1] = 10'b0110010111;
    16'b1000000000010101: out_v[1] = 10'b1100010011;
    16'b1000000000000101: out_v[1] = 10'b0100010111;
    16'b0000000000000010: out_v[1] = 10'b0010001001;
    16'b0100001010010110: out_v[1] = 10'b0111010111;
    16'b1000000010000101: out_v[1] = 10'b1101111111;
    16'b1000000010000110: out_v[1] = 10'b1100110111;
    16'b1000000000010110: out_v[1] = 10'b1100010100;
    16'b1000000000010010: out_v[1] = 10'b0111001111;
    16'b1100000000010110: out_v[1] = 10'b0100010101;
    16'b1000001010010110: out_v[1] = 10'b1010110010;
    16'b1000000000000110: out_v[1] = 10'b0001010101;
    16'b1100000010010110: out_v[1] = 10'b0011011011;
    16'b1000000000011101: out_v[1] = 10'b1101000011;
    16'b0000000000010011: out_v[1] = 10'b1110011110;
    16'b0000000000010001: out_v[1] = 10'b0101001101;
    16'b0000000010010010: out_v[1] = 10'b0101100101;
    16'b1100000010000110: out_v[1] = 10'b1111001110;
    16'b0000000000010010: out_v[1] = 10'b1001001101;
    16'b0000000010000110: out_v[1] = 10'b1100000111;
    16'b1000000010010100: out_v[1] = 10'b1001001001;
    16'b1100001010010110: out_v[1] = 10'b0111010001;
    16'b1100000010010111: out_v[1] = 10'b0011010101;
    16'b1000000000000010: out_v[1] = 10'b0111010111;
    16'b0000000000010110: out_v[1] = 10'b1001111100;
    16'b0000001010000110: out_v[1] = 10'b0111100010;
    16'b0000001010010100: out_v[1] = 10'b0010100011;
    16'b1000000000010100: out_v[1] = 10'b1010010110;
    16'b1000000000010001: out_v[1] = 10'b1111011111;
    16'b0100001010010100: out_v[1] = 10'b1011011110;
    16'b0000000010010100: out_v[1] = 10'b0010110001;
    16'b1000000000010011: out_v[1] = 10'b1110110010;
    16'b1000000010010010: out_v[1] = 10'b0010110001;
    16'b1100000000010111: out_v[1] = 10'b1111100011;
    16'b1100001010010111: out_v[1] = 10'b1010110011;
    16'b0100001000000000: out_v[1] = 10'b0001110011;
    16'b0100000000010000: out_v[1] = 10'b0111011100;
    16'b0000000000010000: out_v[1] = 10'b0000110111;
    16'b0100000000000000: out_v[1] = 10'b1000011110;
    16'b0100001010010000: out_v[1] = 10'b1001010111;
    16'b0000000000000000: out_v[1] = 10'b1001011000;
    16'b0100001000010000: out_v[1] = 10'b1001100111;
    16'b0100000010010000: out_v[1] = 10'b1100010010;
    16'b0000000010010000: out_v[1] = 10'b0011100110;
    16'b0100001000010100: out_v[1] = 10'b1011001000;
    16'b1000001000010110: out_v[1] = 10'b0111010000;
    16'b1100001000000110: out_v[1] = 10'b0000010011;
    16'b0100001000010110: out_v[1] = 10'b1100001011;
    16'b0000001000010010: out_v[1] = 10'b1001100110;
    16'b0000000000010100: out_v[1] = 10'b0010110110;
    16'b0100000000000100: out_v[1] = 10'b1111100010;
    16'b1000001000000100: out_v[1] = 10'b0111101011;
    16'b0100000000010100: out_v[1] = 10'b0110011011;
    16'b0100001000000100: out_v[1] = 10'b0010010110;
    16'b0000001000000110: out_v[1] = 10'b0010110101;
    16'b0000001000000100: out_v[1] = 10'b0101010000;
    16'b1000001000010100: out_v[1] = 10'b0000101100;
    16'b0000001000010100: out_v[1] = 10'b1100001000;
    16'b0000001000010111: out_v[1] = 10'b0101011011;
    16'b0000001000010000: out_v[1] = 10'b0000001100;
    16'b1000001000010111: out_v[1] = 10'b0010110110;
    16'b1000001000000110: out_v[1] = 10'b1011101000;
    16'b1000000000000100: out_v[1] = 10'b1100110110;
    16'b0100001000010010: out_v[1] = 10'b1011100101;
    16'b0100000000010110: out_v[1] = 10'b0010011001;
    16'b1100001000010100: out_v[1] = 10'b0010000100;
    16'b1000001000010010: out_v[1] = 10'b0101100100;
    16'b0000001000000000: out_v[1] = 10'b0110110101;
    16'b0000001000010110: out_v[1] = 10'b1010010100;
    16'b0000001000000010: out_v[1] = 10'b0111000010;
    16'b0100001000000010: out_v[1] = 10'b0110111111;
    16'b1100000000000100: out_v[1] = 10'b0111011010;
    16'b1100001000010110: out_v[1] = 10'b1010100111;
    16'b0100001000000110: out_v[1] = 10'b0100110000;
    16'b0100101000010000: out_v[1] = 10'b0001010101;
    16'b1100000000010100: out_v[1] = 10'b1011000110;
    16'b0000000000000110: out_v[1] = 10'b0000110111;
    16'b1100001010010100: out_v[1] = 10'b1000001001;
    16'b0100000010000100: out_v[1] = 10'b0111100110;
    16'b1000001010010000: out_v[1] = 10'b0111100000;
    16'b1100001010000100: out_v[1] = 10'b1011110110;
    16'b0100000010010100: out_v[1] = 10'b0111110100;
    16'b0100001010000100: out_v[1] = 10'b0000111010;
    16'b1000001010010100: out_v[1] = 10'b0001101000;
    16'b1100001000010000: out_v[1] = 10'b0100011001;
    16'b0000001010000100: out_v[1] = 10'b0000100110;
    16'b1100001010000000: out_v[1] = 10'b1100001111;
    16'b1100001010010000: out_v[1] = 10'b1101000010;
    16'b1000001010000000: out_v[1] = 10'b1010100110;
    16'b1100000010010000: out_v[1] = 10'b0011101000;
    16'b1100000010010100: out_v[1] = 10'b1001111000;
    16'b0100000010000000: out_v[1] = 10'b0110111100;
    16'b1100000010000100: out_v[1] = 10'b1011001100;
    16'b1000001010000100: out_v[1] = 10'b1000101001;
    16'b1100001000000100: out_v[1] = 10'b1110000111;
    16'b0100001010000000: out_v[1] = 10'b0000110001;
    16'b0100001010000110: out_v[1] = 10'b0101110010;
    16'b0100001010000010: out_v[1] = 10'b1100010001;
    16'b0000001010010000: out_v[1] = 10'b1100001000;
    16'b0000001010000010: out_v[1] = 10'b1010101111;
    16'b1100001000000111: out_v[1] = 10'b0000011011;
    16'b0100001010010010: out_v[1] = 10'b0110010110;
    16'b0000001010010010: out_v[1] = 10'b1110011010;
    16'b0000001000000011: out_v[1] = 10'b0111101111;
    16'b1100001010000110: out_v[1] = 10'b0111000011;
    16'b1000001000000111: out_v[1] = 10'b1101101110;
    16'b0000001010000000: out_v[1] = 10'b1100011000;
    16'b0000001010010011: out_v[1] = 10'b0111111100;
    16'b0000001010000011: out_v[1] = 10'b1001110011;
    16'b0100001000000111: out_v[1] = 10'b1010101110;
    16'b0000001000000111: out_v[1] = 10'b0010111111;
    16'b0000001000001111: out_v[1] = 10'b1101011101;
    16'b0100001000000011: out_v[1] = 10'b0101100110;
    16'b0100001010000011: out_v[1] = 10'b1000110011;
    16'b0010000010000000: out_v[1] = 10'b1011011110;
    16'b0100000010000010: out_v[1] = 10'b1000100110;
    16'b0010000010010000: out_v[1] = 10'b1001011011;
    16'b1010001010010100: out_v[1] = 10'b0111111011;
    16'b0110001010010100: out_v[1] = 10'b0111000010;
    16'b0110000010000000: out_v[1] = 10'b1010100110;
    16'b0010001010010100: out_v[1] = 10'b0010010110;
    16'b0000000010000000: out_v[1] = 10'b1001100010;
    16'b0010001010000100: out_v[1] = 10'b0111011111;
    16'b1000001000010000: out_v[1] = 10'b1100001000;
    16'b0010000010010100: out_v[1] = 10'b1010001011;
    16'b0100000000000010: out_v[1] = 10'b1101001010;
    16'b0000000010000100: out_v[1] = 10'b1110001011;
    16'b1000001010010010: out_v[1] = 10'b1011001100;
    16'b1000001010000110: out_v[1] = 10'b1111010000;
    16'b1100000000000110: out_v[1] = 10'b0011001000;
    16'b0001001000000000: out_v[1] = 10'b1001000011;
    16'b0101001010010000: out_v[1] = 10'b0101000011;
    16'b0101001000010100: out_v[1] = 10'b1101101011;
    16'b0101001010000000: out_v[1] = 10'b0111001101;
    16'b0101001000010000: out_v[1] = 10'b0101010011;
    16'b0101001000000000: out_v[1] = 10'b0100100010;
    16'b0101000000010000: out_v[1] = 10'b1011010111;
    16'b0001001000010100: out_v[1] = 10'b1101101101;
    16'b0001001000010000: out_v[1] = 10'b0111011100;
    16'b0101001000000100: out_v[1] = 10'b1001111111;
    16'b0000001100010000: out_v[1] = 10'b0010101011;
    16'b0101001010000100: out_v[1] = 10'b0111100101;
    16'b0001001000000100: out_v[1] = 10'b1001011111;
    16'b0100001010001100: out_v[1] = 10'b0110001011;
    16'b0010001010010000: out_v[1] = 10'b0111000111;
    16'b0110001010010000: out_v[1] = 10'b1001011111;
    16'b0100001000010111: out_v[1] = 10'b1011000011;
    default: out_v[1] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0101000001000000: out_v[2] = 10'b1010110110;
    16'b0100000011000000: out_v[2] = 10'b0010001011;
    16'b0100000010001000: out_v[2] = 10'b0000001100;
    16'b1100000010001000: out_v[2] = 10'b0011111110;
    16'b0100000001000000: out_v[2] = 10'b1010000010;
    16'b0100000000000000: out_v[2] = 10'b1011011001;
    16'b0100000011001000: out_v[2] = 10'b0101000001;
    16'b0000000001000000: out_v[2] = 10'b0100110100;
    16'b0000000010001000: out_v[2] = 10'b0100001101;
    16'b0000000000000000: out_v[2] = 10'b1111000000;
    16'b0000000011001000: out_v[2] = 10'b0000101000;
    16'b0000000011000000: out_v[2] = 10'b0101110011;
    16'b0100000010000000: out_v[2] = 10'b1110000111;
    16'b1100000001000000: out_v[2] = 10'b1011100001;
    16'b1100000011000000: out_v[2] = 10'b1111100110;
    16'b1000000010000000: out_v[2] = 10'b0010001011;
    16'b0000000010000000: out_v[2] = 10'b1011100110;
    16'b1100000000000000: out_v[2] = 10'b1001011011;
    16'b0101000000000000: out_v[2] = 10'b1110111000;
    16'b0001000010000000: out_v[2] = 10'b1010011111;
    16'b1000000000000000: out_v[2] = 10'b1100110110;
    16'b0001000010001000: out_v[2] = 10'b1110000101;
    16'b1100000011001000: out_v[2] = 10'b1000010110;
    16'b0101000011000000: out_v[2] = 10'b0110011011;
    16'b1000000010001000: out_v[2] = 10'b1110100011;
    16'b1100100000000000: out_v[2] = 10'b0011110111;
    16'b1100000010000000: out_v[2] = 10'b0101010010;
    16'b1000000001000000: out_v[2] = 10'b0101000111;
    16'b1000000011001000: out_v[2] = 10'b1011011111;
    16'b1000000011000000: out_v[2] = 10'b1100101100;
    16'b0000100000000000: out_v[2] = 10'b0101010100;
    16'b0001000000000000: out_v[2] = 10'b1110001011;
    16'b1001000000000000: out_v[2] = 10'b1110001101;
    16'b1011100000000000: out_v[2] = 10'b1111111011;
    16'b1000100010000000: out_v[2] = 10'b1100100011;
    16'b1100100010001000: out_v[2] = 10'b1000000100;
    16'b1000100000000000: out_v[2] = 10'b1000001100;
    16'b0011000000000000: out_v[2] = 10'b0101100100;
    16'b1011000010000000: out_v[2] = 10'b1011010101;
    16'b1000100010001000: out_v[2] = 10'b0110100100;
    16'b1001100000000000: out_v[2] = 10'b0110001101;
    16'b0000000000001000: out_v[2] = 10'b1101000011;
    16'b1000100010000001: out_v[2] = 10'b0100101111;
    16'b1100100010000000: out_v[2] = 10'b1011000010;
    16'b0100000000001000: out_v[2] = 10'b0101000111;
    16'b1011100010000000: out_v[2] = 10'b1110110011;
    16'b1000100000000001: out_v[2] = 10'b1001001110;
    16'b0000000000000001: out_v[2] = 10'b1100100111;
    16'b0001000011000000: out_v[2] = 10'b1010011110;
    16'b0001000001000000: out_v[2] = 10'b0110111010;
    16'b1000100011001000: out_v[2] = 10'b1101100101;
    16'b0011000001000000: out_v[2] = 10'b0100111010;
    16'b0011000010000000: out_v[2] = 10'b0010011111;
    16'b1000100011000000: out_v[2] = 10'b1000111110;
    16'b1000100001000000: out_v[2] = 10'b0000001000;
    16'b0111000000000000: out_v[2] = 10'b1011001110;
    16'b0110000000000000: out_v[2] = 10'b1001010010;
    16'b0111000001000000: out_v[2] = 10'b1110100001;
    16'b0010000000000000: out_v[2] = 10'b0100011010;
    16'b0011000011000000: out_v[2] = 10'b1101100010;
    16'b0100100000000000: out_v[2] = 10'b1001101001;
    16'b1100100001000000: out_v[2] = 10'b1100101110;
    16'b0000100001000000: out_v[2] = 10'b1011100011;
    16'b0100100001000000: out_v[2] = 10'b1011000011;
    16'b1001000001000000: out_v[2] = 10'b1011010010;
    default: out_v[2] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0101000010000000: out_v[3] = 10'b1101000011;
    16'b0100010010000000: out_v[3] = 10'b0100000100;
    16'b0001010000000000: out_v[3] = 10'b1000001011;
    16'b0101010000000000: out_v[3] = 10'b1101100001;
    16'b0101000000000000: out_v[3] = 10'b1100100110;
    16'b0001000010000000: out_v[3] = 10'b0100110011;
    16'b0001000000000000: out_v[3] = 10'b0011110100;
    16'b0100010000000000: out_v[3] = 10'b1000101100;
    16'b0101010010000000: out_v[3] = 10'b0011100100;
    16'b0100000010000000: out_v[3] = 10'b1100010111;
    16'b0100000000000000: out_v[3] = 10'b0111011001;
    16'b0000010000000000: out_v[3] = 10'b1000001111;
    16'b0000000000000000: out_v[3] = 10'b0010010110;
    16'b0000000010000000: out_v[3] = 10'b0101101101;
    16'b0000010010000000: out_v[3] = 10'b0111001011;
    16'b0100000000010000: out_v[3] = 10'b1010110100;
    16'b0100010010010000: out_v[3] = 10'b1100001101;
    16'b0110000010010000: out_v[3] = 10'b1011001111;
    16'b0100010000010000: out_v[3] = 10'b1101111011;
    16'b0100000010010000: out_v[3] = 10'b0011001011;
    16'b0110010000010000: out_v[3] = 10'b1010001010;
    16'b0110010010010000: out_v[3] = 10'b0111100110;
    16'b0110000000010000: out_v[3] = 10'b0010101100;
    16'b0010000000010000: out_v[3] = 10'b0011001110;
    16'b1100010000000000: out_v[3] = 10'b1110111011;
    16'b0000000000010000: out_v[3] = 10'b1101000110;
    16'b0000000010010000: out_v[3] = 10'b0001011010;
    16'b0101000000100000: out_v[3] = 10'b0111110110;
    16'b0101010000100000: out_v[3] = 10'b1101011110;
    16'b0010000010010000: out_v[3] = 10'b1111010010;
    16'b0001000000000010: out_v[3] = 10'b1110001000;
    16'b0000000000000010: out_v[3] = 10'b0110011011;
    16'b0001010010000000: out_v[3] = 10'b0111011010;
    default: out_v[3] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000000000001: out_v[4] = 10'b1100000110;
    16'b0010000100000001: out_v[4] = 10'b0011100001;
    16'b0010000101000011: out_v[4] = 10'b0000100001;
    16'b0010000101000001: out_v[4] = 10'b0010110001;
    16'b0010000000000001: out_v[4] = 10'b1010010001;
    16'b0010000001000001: out_v[4] = 10'b1000110001;
    16'b0010000001000011: out_v[4] = 10'b1000011011;
    16'b0000000101000011: out_v[4] = 10'b0000111011;
    16'b0010000000000000: out_v[4] = 10'b0011001110;
    16'b0010000100000000: out_v[4] = 10'b0001111110;
    16'b0000000001000001: out_v[4] = 10'b0010101110;
    16'b0000000001000000: out_v[4] = 10'b1011101011;
    16'b0000000000000000: out_v[4] = 10'b0000110010;
    16'b0010000101000000: out_v[4] = 10'b1111001100;
    16'b0000000101000000: out_v[4] = 10'b0010010111;
    16'b0000000101000001: out_v[4] = 10'b0000011111;
    16'b0010000001000000: out_v[4] = 10'b1100100110;
    16'b0000000100000000: out_v[4] = 10'b1011001011;
    16'b0001001000000000: out_v[4] = 10'b0100001000;
    16'b0011001000000000: out_v[4] = 10'b0111100110;
    16'b0000001000000000: out_v[4] = 10'b0001100101;
    16'b0110000100000000: out_v[4] = 10'b0011111111;
    16'b0001000000000000: out_v[4] = 10'b1010100101;
    16'b0100000100000000: out_v[4] = 10'b0000011000;
    16'b0011001001000000: out_v[4] = 10'b1001000111;
    16'b0001001100000000: out_v[4] = 10'b0010110110;
    16'b0000000100000001: out_v[4] = 10'b0100000110;
    16'b0100000000000000: out_v[4] = 10'b1000001011;
    16'b0001001000000001: out_v[4] = 10'b1011001011;
    16'b0110000000000000: out_v[4] = 10'b1110011010;
    16'b0010001000000001: out_v[4] = 10'b1100011000;
    16'b0011001001000001: out_v[4] = 10'b1001101111;
    16'b0011000001000001: out_v[4] = 10'b1011001111;
    16'b0010001001000001: out_v[4] = 10'b0111011101;
    16'b0011001000000001: out_v[4] = 10'b0011001111;
    16'b0000001000000001: out_v[4] = 10'b1011001110;
    16'b0000000000001000: out_v[4] = 10'b0111111011;
    16'b0011000000000001: out_v[4] = 10'b1011000011;
    16'b0010000000001000: out_v[4] = 10'b1111010010;
    default: out_v[4] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100001000010100: out_v[5] = 10'b1011101011;
    16'b0101001000010010: out_v[5] = 10'b0010100111;
    16'b0100011000010100: out_v[5] = 10'b1011111000;
    16'b0100000000000100: out_v[5] = 10'b0101010001;
    16'b0000001000000100: out_v[5] = 10'b1110100101;
    16'b0100010000000000: out_v[5] = 10'b0111110100;
    16'b0000000000000100: out_v[5] = 10'b0101101111;
    16'b0000000000000000: out_v[5] = 10'b0101101011;
    16'b0101011000010000: out_v[5] = 10'b1111001011;
    16'b0100001000000100: out_v[5] = 10'b0001101000;
    16'b0100011000000000: out_v[5] = 10'b0001010111;
    16'b0100001000010010: out_v[5] = 10'b1000100100;
    16'b0100001000000010: out_v[5] = 10'b0011100011;
    16'b0100000000010000: out_v[5] = 10'b0011100100;
    16'b0100000000010100: out_v[5] = 10'b1001001110;
    16'b0100011000010000: out_v[5] = 10'b1110100100;
    16'b0000001000010100: out_v[5] = 10'b0111001001;
    16'b0101011000010100: out_v[5] = 10'b0010001001;
    16'b0100011000000100: out_v[5] = 10'b0001011110;
    16'b0100010000000100: out_v[5] = 10'b0011110101;
    16'b0100010000010100: out_v[5] = 10'b0011110000;
    16'b0100001000000000: out_v[5] = 10'b1101110010;
    16'b0000000000000010: out_v[5] = 10'b1101001101;
    16'b0000000000010000: out_v[5] = 10'b1110100101;
    16'b0000000000010100: out_v[5] = 10'b0100001100;
    16'b0101001000010110: out_v[5] = 10'b1111100110;
    16'b0101011000000100: out_v[5] = 10'b1001010010;
    16'b0101001000010100: out_v[5] = 10'b0111111111;
    16'b0101000000000010: out_v[5] = 10'b0100011101;
    16'b0101001000000100: out_v[5] = 10'b1011011111;
    16'b0000001000000000: out_v[5] = 10'b1110001100;
    16'b0100001000010110: out_v[5] = 10'b0101000110;
    16'b0100001000010000: out_v[5] = 10'b0110111100;
    16'b0101001000000010: out_v[5] = 10'b0110000001;
    16'b0100000000000000: out_v[5] = 10'b0011111011;
    16'b0000001000000010: out_v[5] = 10'b0110101011;
    16'b0101011000000000: out_v[5] = 10'b0010111111;
    16'b0001011000010100: out_v[5] = 10'b0000010001;
    16'b0000010000000100: out_v[5] = 10'b1001011011;
    16'b0001000000000100: out_v[5] = 10'b0001101111;
    16'b0001010000000100: out_v[5] = 10'b0000110011;
    16'b0000000000000110: out_v[5] = 10'b1111000011;
    16'b0001000000000110: out_v[5] = 10'b0110011001;
    16'b0001000000000000: out_v[5] = 10'b0011011001;
    16'b0100000100000100: out_v[5] = 10'b0001010101;
    16'b0101010000010100: out_v[5] = 10'b0011110100;
    16'b0000010000010100: out_v[5] = 10'b1101001100;
    16'b0000000100000100: out_v[5] = 10'b0001111111;
    16'b0101000000000100: out_v[5] = 10'b1000110100;
    16'b0001010000010100: out_v[5] = 10'b1001110110;
    16'b0101000000010100: out_v[5] = 10'b0101000101;
    16'b0101010000000100: out_v[5] = 10'b1111110111;
    16'b0001000000010100: out_v[5] = 10'b1011100010;
    16'b0100000100010100: out_v[5] = 10'b0000111110;
    16'b0100010000010000: out_v[5] = 10'b0111110110;
    16'b0000011000010100: out_v[5] = 10'b0011000110;
    16'b0101001000000000: out_v[5] = 10'b1111000111;
    16'b0101001000010000: out_v[5] = 10'b1111010001;
    16'b0001000000010010: out_v[5] = 10'b1000101011;
    16'b0100000000000010: out_v[5] = 10'b0001111010;
    16'b0101000000000000: out_v[5] = 10'b0011111011;
    16'b0000001000010010: out_v[5] = 10'b1100001110;
    16'b0000001000010000: out_v[5] = 10'b0101110110;
    16'b0000000000010010: out_v[5] = 10'b1101100011;
    16'b0101000000010010: out_v[5] = 10'b0100011100;
    16'b0100000000010010: out_v[5] = 10'b0000001011;
    16'b0001001000010010: out_v[5] = 10'b0101001001;
    16'b0001000000000010: out_v[5] = 10'b1000110001;
    16'b0101000000010000: out_v[5] = 10'b0011111010;
    16'b0001001000000010: out_v[5] = 10'b0010001011;
    16'b0000001000010110: out_v[5] = 10'b0010111010;
    16'b0000011000000000: out_v[5] = 10'b0111011001;
    16'b0000000100010000: out_v[5] = 10'b1000000010;
    16'b0000000000010110: out_v[5] = 10'b0010000010;
    16'b0000011000010000: out_v[5] = 10'b1100111000;
    16'b0000001000000110: out_v[5] = 10'b1000000111;
    16'b0000010000010000: out_v[5] = 10'b0011111000;
    16'b0100001000000110: out_v[5] = 10'b0110011011;
    16'b0001001000000100: out_v[5] = 10'b1100110110;
    16'b0000011000000100: out_v[5] = 10'b0111010011;
    16'b0100001010010000: out_v[5] = 10'b1111001110;
    16'b0100000010010000: out_v[5] = 10'b1111001100;
    16'b0100001010000000: out_v[5] = 10'b1111001010;
    16'b0100000010000000: out_v[5] = 10'b1011010011;
    16'b0100000000010110: out_v[5] = 10'b0100011111;
    16'b0001000000010110: out_v[5] = 10'b1011100110;
    16'b0100000000110000: out_v[5] = 10'b0111010111;
    16'b0000000010010000: out_v[5] = 10'b1110110011;
    16'b0000000010000000: out_v[5] = 10'b0110111011;
    16'b0001001000010110: out_v[5] = 10'b1101000001;
    16'b0001001000000110: out_v[5] = 10'b0101100110;
    16'b0100000000000110: out_v[5] = 10'b1001110111;
    default: out_v[5] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1011000010110111: out_v[6] = 10'b0100001100;
    16'b1011000010110001: out_v[6] = 10'b0001111111;
    16'b0011001000010001: out_v[6] = 10'b0011011011;
    16'b0011001010010001: out_v[6] = 10'b0011100011;
    16'b0011000010110001: out_v[6] = 10'b1110110110;
    16'b1011001010110101: out_v[6] = 10'b1011110001;
    16'b1010000010110101: out_v[6] = 10'b1011111110;
    16'b1011001010110001: out_v[6] = 10'b1000101111;
    16'b1010001010110001: out_v[6] = 10'b0010001011;
    16'b1001001100110001: out_v[6] = 10'b0110100001;
    16'b1011000010110011: out_v[6] = 10'b0001111001;
    16'b1011000010110101: out_v[6] = 10'b1010110110;
    16'b1011000000110001: out_v[6] = 10'b0110111110;
    16'b1010000010110001: out_v[6] = 10'b1011011111;
    16'b1011001000010001: out_v[6] = 10'b0101000110;
    16'b0011001010000001: out_v[6] = 10'b1110010110;
    16'b0011001100000001: out_v[6] = 10'b1011011110;
    16'b0011000010110011: out_v[6] = 10'b1100001001;
    16'b1001001000110001: out_v[6] = 10'b1000100011;
    16'b1001000000110001: out_v[6] = 10'b0010011001;
    16'b0011001010010101: out_v[6] = 10'b0101110110;
    16'b1011001100110001: out_v[6] = 10'b0111000111;
    16'b0001000010110001: out_v[6] = 10'b1101111101;
    16'b0011001010110001: out_v[6] = 10'b1111101111;
    16'b0010001010010001: out_v[6] = 10'b0110111011;
    16'b0011001000000001: out_v[6] = 10'b1100010001;
    16'b1011001000110101: out_v[6] = 10'b0101100010;
    16'b0010000010110001: out_v[6] = 10'b1110110111;
    16'b0010001010110001: out_v[6] = 10'b1110100110;
    16'b0011001110010001: out_v[6] = 10'b0111011010;
    16'b0011000010110101: out_v[6] = 10'b0001001111;
    16'b0011000000110001: out_v[6] = 10'b1001110101;
    16'b1011001000110001: out_v[6] = 10'b0001110101;
    16'b0011001110110001: out_v[6] = 10'b1101100011;
    16'b1010000000110001: out_v[6] = 10'b1111001010;
    16'b1011001010010001: out_v[6] = 10'b1100011111;
    16'b1011000010100001: out_v[6] = 10'b0111000111;
    16'b1011000000110101: out_v[6] = 10'b1000011110;
    16'b0011001110000001: out_v[6] = 10'b1110110101;
    16'b1001001100000001: out_v[6] = 10'b1011011001;
    16'b0011000100000001: out_v[6] = 10'b0001100011;
    16'b0011000100000101: out_v[6] = 10'b0101001101;
    16'b0000000000000000: out_v[6] = 10'b1001011110;
    16'b1000000000000000: out_v[6] = 10'b0010001111;
    16'b0001000000000001: out_v[6] = 10'b1111000111;
    16'b0001000100000100: out_v[6] = 10'b1100100011;
    16'b0000000100000000: out_v[6] = 10'b1011001100;
    16'b0001000000000000: out_v[6] = 10'b1101000001;
    16'b0001000100000000: out_v[6] = 10'b1100100001;
    16'b0000000000000100: out_v[6] = 10'b0100110011;
    16'b0001000100000101: out_v[6] = 10'b0011011001;
    16'b1001000000000000: out_v[6] = 10'b0000101101;
    16'b0011000110000001: out_v[6] = 10'b1111000010;
    16'b0001000100000001: out_v[6] = 10'b0010011010;
    16'b0001000000000100: out_v[6] = 10'b1110101000;
    16'b1000000100000000: out_v[6] = 10'b1001011100;
    16'b0011000100000000: out_v[6] = 10'b1110110111;
    16'b0001000000000101: out_v[6] = 10'b0011110101;
    16'b0011000000000001: out_v[6] = 10'b1001011011;
    16'b1001000100000000: out_v[6] = 10'b0000111011;
    16'b0011001010100001: out_v[6] = 10'b0111011001;
    16'b1011000100000001: out_v[6] = 10'b0000100101;
    16'b0001001100000001: out_v[6] = 10'b1010100001;
    16'b0011000110100001: out_v[6] = 10'b1011000111;
    16'b0010001010000001: out_v[6] = 10'b1110101011;
    16'b0011001100100001: out_v[6] = 10'b1110101100;
    16'b1011000110000001: out_v[6] = 10'b0000111110;
    16'b0010000110000001: out_v[6] = 10'b1101111011;
    16'b1001000100000001: out_v[6] = 10'b0011001100;
    16'b0010001110000001: out_v[6] = 10'b0100001011;
    16'b0011001110100001: out_v[6] = 10'b0001101010;
    16'b0001000110100001: out_v[6] = 10'b1000110111;
    16'b0000000100100000: out_v[6] = 10'b1100000111;
    16'b0000001110000001: out_v[6] = 10'b0111011110;
    16'b0001001110100001: out_v[6] = 10'b0001011010;
    16'b0001000110000001: out_v[6] = 10'b0011100101;
    16'b0010001110000000: out_v[6] = 10'b0110111100;
    16'b0010001100000000: out_v[6] = 10'b1101000111;
    16'b0001000100100000: out_v[6] = 10'b1111001001;
    16'b0010000100000000: out_v[6] = 10'b1100000101;
    16'b0011000010000001: out_v[6] = 10'b0001011111;
    16'b0001001110000001: out_v[6] = 10'b0111110110;
    16'b1010000110000001: out_v[6] = 10'b1001110111;
    16'b0011000100100001: out_v[6] = 10'b1010110111;
    16'b0000001110000000: out_v[6] = 10'b1110110011;
    16'b0000000110000001: out_v[6] = 10'b1010101111;
    16'b0010000100000001: out_v[6] = 10'b1100011101;
    16'b0010001100000001: out_v[6] = 10'b1011011101;
    16'b0010001110100001: out_v[6] = 10'b1001100100;
    16'b0011000100100000: out_v[6] = 10'b1011110010;
    16'b1011001110000001: out_v[6] = 10'b1010101110;
    16'b0001000110100000: out_v[6] = 10'b0101111010;
    16'b0001000100100001: out_v[6] = 10'b0100000100;
    16'b1011001000000101: out_v[6] = 10'b1010100101;
    16'b1011000000000000: out_v[6] = 10'b1111110010;
    16'b1001000100000101: out_v[6] = 10'b0000111011;
    16'b1011001010100001: out_v[6] = 10'b0010001000;
    16'b1011000000000101: out_v[6] = 10'b1011010111;
    16'b0010001000000001: out_v[6] = 10'b0000100011;
    16'b0010000000000001: out_v[6] = 10'b1101010001;
    16'b1011000000000100: out_v[6] = 10'b1111011101;
    16'b0010000010000001: out_v[6] = 10'b1000011010;
    16'b1000001000100000: out_v[6] = 10'b0000111010;
    16'b1001000000000100: out_v[6] = 10'b1001011101;
    16'b1011001000010101: out_v[6] = 10'b0101100011;
    16'b1011000100000101: out_v[6] = 10'b1010010101;
    16'b1011001010100101: out_v[6] = 10'b1000010001;
    16'b1011001000100001: out_v[6] = 10'b0100011010;
    16'b0011000000000101: out_v[6] = 10'b0011011111;
    16'b1011000010000101: out_v[6] = 10'b1111011010;
    16'b1011001000100101: out_v[6] = 10'b0011110110;
    16'b1011001000100000: out_v[6] = 10'b0111011011;
    16'b1011000010000001: out_v[6] = 10'b0001011101;
    16'b1011000000000001: out_v[6] = 10'b1010101010;
    16'b1001000000000101: out_v[6] = 10'b0101111000;
    16'b1010001000100000: out_v[6] = 10'b1101100011;
    16'b0011001000100001: out_v[6] = 10'b0011011111;
    16'b0010000000000000: out_v[6] = 10'b0000110011;
    16'b0010000000000101: out_v[6] = 10'b1010101111;
    16'b1010001000000000: out_v[6] = 10'b1011110110;
    16'b1011001010000001: out_v[6] = 10'b0011000110;
    16'b1011001010000101: out_v[6] = 10'b0011111110;
    16'b1011001000000001: out_v[6] = 10'b0101010111;
    16'b0011001000000101: out_v[6] = 10'b1111110100;
    16'b1010000000000101: out_v[6] = 10'b1010011110;
    16'b1011000000010101: out_v[6] = 10'b1011011000;
    16'b1000000000000100: out_v[6] = 10'b0111101100;
    16'b1011000000100101: out_v[6] = 10'b1110100011;
    16'b1001001100010001: out_v[6] = 10'b1000101111;
    16'b0001001100010101: out_v[6] = 10'b1100101110;
    16'b0001000100110001: out_v[6] = 10'b0100111011;
    16'b0000000000010100: out_v[6] = 10'b1011011011;
    16'b0001001000010001: out_v[6] = 10'b0100011000;
    16'b0000001100000000: out_v[6] = 10'b1011000110;
    16'b0001001000010101: out_v[6] = 10'b1111001110;
    16'b0001000000010001: out_v[6] = 10'b1011110111;
    16'b0000001000010100: out_v[6] = 10'b0110011001;
    16'b0010001000010100: out_v[6] = 10'b0011011101;
    16'b0001001100110001: out_v[6] = 10'b0000111010;
    16'b1000001000010001: out_v[6] = 10'b1000001101;
    16'b0010001100010100: out_v[6] = 10'b0001111101;
    16'b0001001100010001: out_v[6] = 10'b1100111011;
    16'b1000001100010001: out_v[6] = 10'b1011001111;
    16'b0010000100010000: out_v[6] = 10'b1101010110;
    16'b1001000000010001: out_v[6] = 10'b1101010010;
    16'b0000000100010000: out_v[6] = 10'b1110001110;
    16'b0000000100010001: out_v[6] = 10'b1101101111;
    16'b0000001100110000: out_v[6] = 10'b0011101010;
    16'b0000001000010000: out_v[6] = 10'b0011011000;
    16'b1000001100010000: out_v[6] = 10'b0110011011;
    16'b1000001000010000: out_v[6] = 10'b0110111111;
    16'b1001000100110001: out_v[6] = 10'b1111010010;
    16'b1001000100010001: out_v[6] = 10'b1111001010;
    16'b1001001000010001: out_v[6] = 10'b0110011001;
    16'b0000001100010000: out_v[6] = 10'b0010111010;
    16'b1001001100010000: out_v[6] = 10'b0000011110;
    16'b1001000000010000: out_v[6] = 10'b1100010001;
    16'b0001000100010001: out_v[6] = 10'b1100100111;
    16'b0001001100010000: out_v[6] = 10'b1001101111;
    16'b0000001100010001: out_v[6] = 10'b1000001011;
    16'b0000001000010001: out_v[6] = 10'b0100010101;
    16'b0000000100010100: out_v[6] = 10'b0001011111;
    16'b0000001100110001: out_v[6] = 10'b1111110110;
    16'b0000000000010000: out_v[6] = 10'b0011010100;
    16'b0000001100010100: out_v[6] = 10'b0001111100;
    16'b0010001000010000: out_v[6] = 10'b1010110111;
    16'b0001001000010000: out_v[6] = 10'b1101011010;
    16'b0000001000010101: out_v[6] = 10'b1100111111;
    16'b0000000000010001: out_v[6] = 10'b1001110100;
    16'b0010001100010000: out_v[6] = 10'b0010111100;
    16'b0001001000000001: out_v[6] = 10'b0110111100;
    16'b1011000010010101: out_v[6] = 10'b1001111110;
    16'b0011000000010001: out_v[6] = 10'b0111001111;
    16'b0011000000010101: out_v[6] = 10'b0001001011;
    16'b1011000100010101: out_v[6] = 10'b0010101000;
    16'b1001000100010101: out_v[6] = 10'b0001010101;
    16'b1011000010010001: out_v[6] = 10'b0100010000;
    16'b0011000010010001: out_v[6] = 10'b0000111010;
    16'b0011000100010101: out_v[6] = 10'b0111100011;
    16'b0000000010000000: out_v[6] = 10'b1111010010;
    16'b0001000010000001: out_v[6] = 10'b1010100010;
    16'b0011000010000000: out_v[6] = 10'b1010111001;
    16'b0010001000000000: out_v[6] = 10'b0011110000;
    16'b0011000010000101: out_v[6] = 10'b1011111001;
    16'b1010001000110001: out_v[6] = 10'b1011011011;
    16'b1000001000110000: out_v[6] = 10'b0111001011;
    16'b1010001010110000: out_v[6] = 10'b1110001110;
    16'b1010001000110000: out_v[6] = 10'b1000100100;
    16'b0001000010000000: out_v[6] = 10'b1111010101;
    16'b1001000000010101: out_v[6] = 10'b0101001110;
    16'b1010000000010101: out_v[6] = 10'b0111010000;
    16'b1010000000000001: out_v[6] = 10'b1010110101;
    16'b0011000010010000: out_v[6] = 10'b1100001011;
    16'b1011000000010001: out_v[6] = 10'b1011011010;
    16'b1000001100000000: out_v[6] = 10'b1001011100;
    16'b0000001100100000: out_v[6] = 10'b1100101101;
    16'b0000000000110000: out_v[6] = 10'b0011011000;
    16'b1000001100110000: out_v[6] = 10'b0011101111;
    16'b0000001000110000: out_v[6] = 10'b0111001000;
    16'b1000000100110000: out_v[6] = 10'b1011111010;
    16'b0000001010110000: out_v[6] = 10'b1111001000;
    16'b1000001100100000: out_v[6] = 10'b1111000011;
    16'b0000001000000000: out_v[6] = 10'b0111100011;
    16'b0000000100110000: out_v[6] = 10'b0101111111;
    16'b0000001110110000: out_v[6] = 10'b1011011010;
    16'b0010001100110000: out_v[6] = 10'b1100111011;
    16'b0000000000100000: out_v[6] = 10'b0001001111;
    16'b0000001000100000: out_v[6] = 10'b0001111110;
    16'b0011001000010101: out_v[6] = 10'b1001001101;
    16'b0001001000000101: out_v[6] = 10'b0000010110;
    16'b1001101000000001: out_v[6] = 10'b1111101011;
    16'b0001000000010101: out_v[6] = 10'b0011110010;
    16'b1001001000000000: out_v[6] = 10'b0110000011;
    16'b0001001000010100: out_v[6] = 10'b0111101111;
    16'b1001001000000001: out_v[6] = 10'b0100010100;
    16'b0011001000000100: out_v[6] = 10'b1101111011;
    16'b0011001100000101: out_v[6] = 10'b1011001111;
    16'b0001001000000000: out_v[6] = 10'b0101110101;
    16'b1001000000000001: out_v[6] = 10'b1110110001;
    16'b0000001000000100: out_v[6] = 10'b1010001101;
    16'b0001001000000100: out_v[6] = 10'b1111100011;
    16'b0001101000000000: out_v[6] = 10'b1101011111;
    16'b1000001000000000: out_v[6] = 10'b0010110001;
    16'b1001101000000000: out_v[6] = 10'b1001111001;
    16'b1001001000010000: out_v[6] = 10'b0111000111;
    16'b0001000000010000: out_v[6] = 10'b0111111010;
    16'b0001101000000101: out_v[6] = 10'b0001111111;
    16'b0001001100000101: out_v[6] = 10'b0010100000;
    16'b0001000000010100: out_v[6] = 10'b1111000111;
    16'b1011000110000101: out_v[6] = 10'b1011000101;
    16'b1000000100000001: out_v[6] = 10'b1110111101;
    16'b1010000100000001: out_v[6] = 10'b1000111011;
    16'b0000000100000101: out_v[6] = 10'b0101000000;
    16'b0011001110000101: out_v[6] = 10'b0101001011;
    16'b1011001110000101: out_v[6] = 10'b0111100010;
    16'b1010000100000101: out_v[6] = 10'b1001110101;
    16'b0010000110000101: out_v[6] = 10'b1110010111;
    16'b0010000110000000: out_v[6] = 10'b1111000011;
    16'b0011000110000101: out_v[6] = 10'b1000111000;
    16'b0010000100000100: out_v[6] = 10'b0100111011;
    16'b0010000100000101: out_v[6] = 10'b1111110001;
    16'b1011001100010101: out_v[6] = 10'b0111000011;
    16'b1010000100000000: out_v[6] = 10'b1011101110;
    16'b1011001100000101: out_v[6] = 10'b1001111001;
    16'b1010000100010101: out_v[6] = 10'b1111100110;
    16'b0001000100010000: out_v[6] = 10'b0010100000;
    16'b1000000000010000: out_v[6] = 10'b1000100010;
    16'b0000000000000101: out_v[6] = 10'b1001100100;
    16'b1001000100010000: out_v[6] = 10'b1101100001;
    16'b0001000100010101: out_v[6] = 10'b1001001100;
    16'b0011001100010101: out_v[6] = 10'b1111000010;
    default: out_v[6] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010000000010001: out_v[7] = 10'b0001100101;
    16'b0110000000010011: out_v[7] = 10'b1000011001;
    16'b0011000100010011: out_v[7] = 10'b1100001111;
    16'b0000000000010011: out_v[7] = 10'b0100000101;
    16'b0010000000000001: out_v[7] = 10'b0110100001;
    16'b0111000100010010: out_v[7] = 10'b0000011101;
    16'b0110000100000011: out_v[7] = 10'b1001011011;
    16'b0110000000000001: out_v[7] = 10'b0000110101;
    16'b0110000100010011: out_v[7] = 10'b1111100110;
    16'b0110000000010001: out_v[7] = 10'b0001001100;
    16'b0010000100010011: out_v[7] = 10'b0110111111;
    16'b0100000100010011: out_v[7] = 10'b0010011111;
    16'b0000000100010010: out_v[7] = 10'b0001011010;
    16'b0110000000000011: out_v[7] = 10'b1101011110;
    16'b0111000100010011: out_v[7] = 10'b0101001000;
    16'b0000000100010011: out_v[7] = 10'b0000101011;
    16'b0010000000000011: out_v[7] = 10'b1010001111;
    16'b0011000100010001: out_v[7] = 10'b0010110011;
    16'b0001000100010001: out_v[7] = 10'b1010011000;
    16'b0111000100010001: out_v[7] = 10'b1001001011;
    16'b0111000100000011: out_v[7] = 10'b1101100000;
    16'b0010000100000011: out_v[7] = 10'b1010000011;
    16'b0010000000010011: out_v[7] = 10'b1010000111;
    16'b0001000100010011: out_v[7] = 10'b0110110011;
    16'b0100000000000011: out_v[7] = 10'b0110001001;
    16'b0100000000010011: out_v[7] = 10'b0111101110;
    16'b0101000100010010: out_v[7] = 10'b0110101111;
    16'b0010000100010001: out_v[7] = 10'b1010100111;
    16'b0111100100010011: out_v[7] = 10'b1000000101;
    16'b0000000100000011: out_v[7] = 10'b0100011011;
    16'b0110000100010010: out_v[7] = 10'b0110011011;
    16'b0000000000000001: out_v[7] = 10'b1010000111;
    16'b0110000000010000: out_v[7] = 10'b0000011111;
    16'b0110000000010010: out_v[7] = 10'b0010011110;
    16'b0010000100010010: out_v[7] = 10'b1001111010;
    16'b0000000000010001: out_v[7] = 10'b0011110101;
    16'b0110100000000001: out_v[7] = 10'b1001100010;
    16'b0110100100010011: out_v[7] = 10'b1000000001;
    16'b0110000100010001: out_v[7] = 10'b1010111011;
    16'b0100100000000001: out_v[7] = 10'b0110010010;
    16'b0110100000000000: out_v[7] = 10'b1100000111;
    16'b0000000000000000: out_v[7] = 10'b0001110110;
    16'b0010000000000000: out_v[7] = 10'b0101001110;
    16'b0110000000000000: out_v[7] = 10'b1100000101;
    16'b0100000000000001: out_v[7] = 10'b0011011010;
    16'b0000100000000000: out_v[7] = 10'b0001110010;
    16'b0010100000000000: out_v[7] = 10'b0101011100;
    16'b0100100001000001: out_v[7] = 10'b0011000111;
    16'b0100000000000000: out_v[7] = 10'b0011100100;
    16'b0100100000000000: out_v[7] = 10'b0110110001;
    16'b0110100000010000: out_v[7] = 10'b1110011010;
    16'b0000100000000001: out_v[7] = 10'b1100110100;
    16'b0100000000010001: out_v[7] = 10'b1111001110;
    16'b0100100000010001: out_v[7] = 10'b1100011110;
    16'b0110100000010001: out_v[7] = 10'b1110100000;
    16'b0100100000010000: out_v[7] = 10'b0100111001;
    16'b0000100000010001: out_v[7] = 10'b1101001110;
    16'b0000000000000011: out_v[7] = 10'b0111000110;
    16'b0000000000010010: out_v[7] = 10'b0101110100;
    16'b0000000000010000: out_v[7] = 10'b1011110010;
    16'b0010100000010001: out_v[7] = 10'b0000100000;
    16'b0000000000000010: out_v[7] = 10'b1000100110;
    16'b0000100000000011: out_v[7] = 10'b0100110110;
    16'b0010100000000001: out_v[7] = 10'b1010001000;
    16'b0100000000010000: out_v[7] = 10'b0110100011;
    16'b0000100000010000: out_v[7] = 10'b1001100110;
    16'b0110100100010000: out_v[7] = 10'b1110011111;
    16'b0110100000010011: out_v[7] = 10'b0110001011;
    16'b0100100100010001: out_v[7] = 10'b1101001000;
    16'b0100100000010011: out_v[7] = 10'b0011011001;
    16'b0110100100010001: out_v[7] = 10'b0110011110;
    16'b0110100000010010: out_v[7] = 10'b1010111110;
    16'b0010100000010000: out_v[7] = 10'b0011011000;
    16'b0010100000010011: out_v[7] = 10'b0100111110;
    16'b0000100100000001: out_v[7] = 10'b0101101001;
    16'b0101100100000001: out_v[7] = 10'b0110110010;
    16'b0000100100000000: out_v[7] = 10'b0001010101;
    16'b0100100100000001: out_v[7] = 10'b0110011000;
    16'b0000100100000010: out_v[7] = 10'b0011010001;
    16'b0101100100010001: out_v[7] = 10'b0111111100;
    16'b0100100100000011: out_v[7] = 10'b0000111011;
    16'b0100100100000000: out_v[7] = 10'b1110000001;
    16'b0001100100000000: out_v[7] = 10'b0001100011;
    16'b0000100001000000: out_v[7] = 10'b1110001000;
    16'b0000100000000010: out_v[7] = 10'b0011100110;
    16'b0001100100000010: out_v[7] = 10'b0011110011;
    16'b0001100100010010: out_v[7] = 10'b0111011000;
    16'b0001100100000001: out_v[7] = 10'b1101011110;
    16'b0000000100010001: out_v[7] = 10'b0011011111;
    16'b0110100100000000: out_v[7] = 10'b0110010101;
    16'b0000000100000000: out_v[7] = 10'b0010011011;
    16'b0001100100010001: out_v[7] = 10'b0110010010;
    16'b0000100100010001: out_v[7] = 10'b1011010101;
    16'b0100100000000011: out_v[7] = 10'b0001011010;
    16'b0001000100010010: out_v[7] = 10'b0100011001;
    16'b0000100100000011: out_v[7] = 10'b1111010010;
    16'b0000000100000010: out_v[7] = 10'b1001111011;
    16'b0001000100000010: out_v[7] = 10'b1101010010;
    16'b0011100100010001: out_v[7] = 10'b0001001111;
    16'b0100000100000000: out_v[7] = 10'b0011101110;
    16'b0010000100000001: out_v[7] = 10'b1111000100;
    16'b0010100100010001: out_v[7] = 10'b0100101110;
    16'b0110000100000001: out_v[7] = 10'b0110010011;
    16'b0100000100000001: out_v[7] = 10'b0011010011;
    16'b0000100100010000: out_v[7] = 10'b1011001011;
    16'b0111100100010001: out_v[7] = 10'b0111110001;
    16'b0010100001010001: out_v[7] = 10'b1110110001;
    16'b0010100000010010: out_v[7] = 10'b0110011010;
    16'b0000100000010010: out_v[7] = 10'b0111100001;
    16'b0000000100010000: out_v[7] = 10'b0011101000;
    16'b0010000000010010: out_v[7] = 10'b1011111110;
    16'b0010000000010000: out_v[7] = 10'b0110001010;
    16'b0000100100010010: out_v[7] = 10'b1011000000;
    16'b0100000001000001: out_v[7] = 10'b1011001010;
    16'b0010100000000010: out_v[7] = 10'b0101011010;
    16'b0010100100010010: out_v[7] = 10'b1011100000;
    16'b0110100000000010: out_v[7] = 10'b0010100100;
    16'b0101100100000011: out_v[7] = 10'b0011011101;
    16'b0100000000000010: out_v[7] = 10'b0000100001;
    16'b0111100100000001: out_v[7] = 10'b0110110010;
    16'b0101100100000000: out_v[7] = 10'b1101100100;
    16'b0110100000000011: out_v[7] = 10'b0010111000;
    16'b0101100000000001: out_v[7] = 10'b0111010011;
    16'b0100000100000010: out_v[7] = 10'b1110000110;
    16'b0101000000000010: out_v[7] = 10'b0110111011;
    16'b0111100000000001: out_v[7] = 10'b1011110111;
    16'b0110100100000001: out_v[7] = 10'b1011101000;
    16'b0101000100000010: out_v[7] = 10'b0010010111;
    16'b0101000000000000: out_v[7] = 10'b1100001010;
    16'b0101000100000000: out_v[7] = 10'b1101100011;
    16'b0111100000000000: out_v[7] = 10'b1001111101;
    16'b0101100100000010: out_v[7] = 10'b0011111110;
    16'b0101100000000000: out_v[7] = 10'b0001100110;
    16'b0010100000000011: out_v[7] = 10'b0111010011;
    16'b0010100100000001: out_v[7] = 10'b1100100110;
    16'b0111100100010000: out_v[7] = 10'b1110010010;
    16'b0110100010000000: out_v[7] = 10'b1001100101;
    16'b0111100110010001: out_v[7] = 10'b1101000001;
    16'b0010100100000011: out_v[7] = 10'b1011100110;
    16'b0011100100000001: out_v[7] = 10'b1011100010;
    16'b0110100100000011: out_v[7] = 10'b1011001111;
    16'b0111100110010000: out_v[7] = 10'b0011000111;
    16'b0111100100000011: out_v[7] = 10'b1100110100;
    16'b0011100100000011: out_v[7] = 10'b1100110010;
    16'b0111100100000000: out_v[7] = 10'b0110010101;
    16'b0101100110010000: out_v[7] = 10'b1101000001;
    16'b0110100110010000: out_v[7] = 10'b1101100111;
    default: out_v[7] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000001000010000: out_v[8] = 10'b0011111100;
    16'b0000001000010010: out_v[8] = 10'b1000111011;
    16'b0000001100010010: out_v[8] = 10'b0110000011;
    16'b0000001100000010: out_v[8] = 10'b1000111000;
    16'b0000001000000010: out_v[8] = 10'b0011111011;
    16'b0000001000000000: out_v[8] = 10'b1111001011;
    16'b0000001100010000: out_v[8] = 10'b0010001111;
    16'b0000000000000110: out_v[8] = 10'b1011001111;
    16'b0000001000010011: out_v[8] = 10'b0111100011;
    16'b0000001100010011: out_v[8] = 10'b0010101011;
    16'b0000001100010110: out_v[8] = 10'b0010111011;
    16'b0000001000000110: out_v[8] = 10'b0110010011;
    16'b0000000000000010: out_v[8] = 10'b1110101001;
    16'b0000001100000110: out_v[8] = 10'b0001011001;
    16'b0000001100000000: out_v[8] = 10'b0001110110;
    16'b0000000100000110: out_v[8] = 10'b1100001011;
    16'b0000000000010010: out_v[8] = 10'b1000111001;
    16'b0000101000010010: out_v[8] = 10'b1100110110;
    16'b0000001100000100: out_v[8] = 10'b1011000110;
    16'b0000101000010000: out_v[8] = 10'b1011010011;
    16'b0000000100001110: out_v[8] = 10'b0010001001;
    16'b0000000100000010: out_v[8] = 10'b0011011111;
    16'b0000000100010110: out_v[8] = 10'b1011110110;
    16'b0000000000000000: out_v[8] = 10'b1001010110;
    16'b0000000000010011: out_v[8] = 10'b0110010000;
    16'b0000000100000100: out_v[8] = 10'b1100101101;
    16'b0000001100001110: out_v[8] = 10'b1010011001;
    16'b0000000100010010: out_v[8] = 10'b0110000011;
    16'b0000000000010000: out_v[8] = 10'b0101101110;
    16'b0000001000010001: out_v[8] = 10'b1001110001;
    16'b0000101000010011: out_v[8] = 10'b1110110011;
    16'b0000000100000000: out_v[8] = 10'b0000001111;
    16'b0000000000000001: out_v[8] = 10'b1111011101;
    16'b0000000000010001: out_v[8] = 10'b1000110010;
    16'b0000000000000011: out_v[8] = 10'b0011001110;
    16'b0000000000001100: out_v[8] = 10'b1000010110;
    16'b0000001000000111: out_v[8] = 10'b0000111110;
    16'b0000001000000100: out_v[8] = 10'b0001101101;
    16'b0000001000001010: out_v[8] = 10'b1011001111;
    16'b0000000000000101: out_v[8] = 10'b0001111001;
    16'b0000000100001100: out_v[8] = 10'b0100110111;
    16'b0000001000001011: out_v[8] = 10'b1011000110;
    16'b0000001000000001: out_v[8] = 10'b0110001100;
    16'b0000001000001100: out_v[8] = 10'b1111010110;
    16'b0000001000000011: out_v[8] = 10'b0010001100;
    16'b0000001000001111: out_v[8] = 10'b1000011111;
    16'b0000101000000010: out_v[8] = 10'b0010110011;
    16'b0000000000001111: out_v[8] = 10'b1001101110;
    16'b0000001000001110: out_v[8] = 10'b1110000110;
    16'b0000001000000101: out_v[8] = 10'b0011111100;
    16'b0000000000000100: out_v[8] = 10'b0010110101;
    16'b0000001100001100: out_v[8] = 10'b0010111101;
    16'b0000001000011111: out_v[8] = 10'b1000101110;
    16'b0000001100000011: out_v[8] = 10'b0101011110;
    16'b0000001000010111: out_v[8] = 10'b0110010000;
    16'b0000100000000010: out_v[8] = 10'b0111010100;
    16'b0000000000000111: out_v[8] = 10'b0000110101;
    16'b0000000000001101: out_v[8] = 10'b0011001011;
    16'b0000000000001110: out_v[8] = 10'b0111100011;
    16'b0000001100001111: out_v[8] = 10'b0000101110;
    16'b0000001100000111: out_v[8] = 10'b1010100011;
    16'b0000101000000001: out_v[8] = 10'b0111001000;
    16'b0000101000000011: out_v[8] = 10'b1111011010;
    16'b0000101000000110: out_v[8] = 10'b1111011110;
    16'b0000001100000001: out_v[8] = 10'b1101001010;
    16'b0000000000011100: out_v[8] = 10'b0001001100;
    16'b0000001000001101: out_v[8] = 10'b0010111011;
    16'b0000001000011101: out_v[8] = 10'b0011001000;
    16'b0010001000000001: out_v[8] = 10'b0001001101;
    16'b0000001100001101: out_v[8] = 10'b1111100001;
    16'b0000101000000101: out_v[8] = 10'b1000110110;
    16'b0000001000010101: out_v[8] = 10'b0110000011;
    16'b0000101000010101: out_v[8] = 10'b1110010111;
    16'b0000001100011101: out_v[8] = 10'b1100010110;
    16'b0000101000010001: out_v[8] = 10'b1110011010;
    16'b0000001000001001: out_v[8] = 10'b0000110110;
    16'b0000001000010100: out_v[8] = 10'b0111001110;
    16'b0000101000001101: out_v[8] = 10'b1110111011;
    16'b0000000000011101: out_v[8] = 10'b0010001001;
    16'b0000001000011100: out_v[8] = 10'b0011100101;
    16'b0000001000010110: out_v[8] = 10'b1010001100;
    16'b0000001100000101: out_v[8] = 10'b0101100000;
    16'b0000100000000001: out_v[8] = 10'b1000001011;
    16'b0000000000011110: out_v[8] = 10'b1110001010;
    16'b0000001100001000: out_v[8] = 10'b0011011010;
    16'b0010000000000001: out_v[8] = 10'b1001011101;
    16'b0000000100000001: out_v[8] = 10'b1000111100;
    16'b0000000100001001: out_v[8] = 10'b1000110011;
    16'b0010000000010001: out_v[8] = 10'b1101110101;
    16'b0000001100001001: out_v[8] = 10'b0100010001;
    16'b0000001100001010: out_v[8] = 10'b0101010010;
    16'b0000000100000101: out_v[8] = 10'b1110000100;
    16'b0010001000010001: out_v[8] = 10'b1011100110;
    16'b0000001100010001: out_v[8] = 10'b1100001101;
    16'b0000000100001101: out_v[8] = 10'b0111100010;
    16'b0000000100000111: out_v[8] = 10'b1111010110;
    16'b0010000000000100: out_v[8] = 10'b0010110101;
    16'b1010001100010000: out_v[8] = 10'b0111111000;
    16'b1010000100010000: out_v[8] = 10'b0101011010;
    16'b0010000100000000: out_v[8] = 10'b0001101011;
    16'b1010000000010000: out_v[8] = 10'b0010000101;
    16'b0000000100010000: out_v[8] = 10'b0011100011;
    16'b0010000000010000: out_v[8] = 10'b0011101111;
    16'b0010001100010000: out_v[8] = 10'b0111110100;
    16'b1010000000000000: out_v[8] = 10'b1001101111;
    16'b0010000100010000: out_v[8] = 10'b1011110011;
    16'b0010000000001100: out_v[8] = 10'b0000110110;
    16'b0010000000000000: out_v[8] = 10'b0111011000;
    16'b1010000100000000: out_v[8] = 10'b0010111111;
    16'b0000001110010000: out_v[8] = 10'b0110111111;
    16'b1000000100010000: out_v[8] = 10'b0110011001;
    16'b0000001101010000: out_v[8] = 10'b0111000101;
    16'b0000000100000011: out_v[8] = 10'b0110100110;
    16'b0000000100001111: out_v[8] = 10'b1100010010;
    16'b0010000000010011: out_v[8] = 10'b0101011111;
    16'b1010000000010001: out_v[8] = 10'b1001000110;
    16'b0010000100000001: out_v[8] = 10'b1100001001;
    16'b1010000000000001: out_v[8] = 10'b1000110111;
    16'b0010001100000001: out_v[8] = 10'b1100001111;
    default: out_v[8] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000000000000: out_v[9] = 10'b1010010010;
    16'b1001000000000000: out_v[9] = 10'b0001111001;
    16'b1001100100100000: out_v[9] = 10'b0111110011;
    16'b1001100000100000: out_v[9] = 10'b0111000001;
    16'b1000000000000000: out_v[9] = 10'b0011100001;
    16'b1001000100000000: out_v[9] = 10'b0010000111;
    16'b1001100100000000: out_v[9] = 10'b1111110100;
    16'b1001000100100000: out_v[9] = 10'b0001011011;
    16'b1001101000100000: out_v[9] = 10'b1011011110;
    16'b0001100000000000: out_v[9] = 10'b1000101110;
    16'b0000101000100000: out_v[9] = 10'b0100010001;
    16'b1001101100100000: out_v[9] = 10'b0101101010;
    16'b1000001000000000: out_v[9] = 10'b0001101001;
    16'b1000001000100000: out_v[9] = 10'b0110101011;
    16'b0000100000100000: out_v[9] = 10'b1100010101;
    16'b1001101000000000: out_v[9] = 10'b0100000110;
    16'b0001100001100000: out_v[9] = 10'b1100110001;
    16'b0000101000000000: out_v[9] = 10'b1000111101;
    16'b1000101000100000: out_v[9] = 10'b0001110101;
    16'b1001000000100000: out_v[9] = 10'b0100011111;
    16'b0000101001100000: out_v[9] = 10'b0111110000;
    16'b1000100000100000: out_v[9] = 10'b0001110110;
    16'b0001100100100000: out_v[9] = 10'b0111011011;
    16'b1001001000000000: out_v[9] = 10'b1101100010;
    16'b1000100100100000: out_v[9] = 10'b0011100111;
    16'b1000000000100000: out_v[9] = 10'b1010010000;
    16'b1001100000000000: out_v[9] = 10'b0110110010;
    16'b0001100000100000: out_v[9] = 10'b0110110100;
    16'b0001101000100000: out_v[9] = 10'b0011111011;
    16'b0000100000000000: out_v[9] = 10'b0001011111;
    16'b0001000000000000: out_v[9] = 10'b0101111011;
    16'b1001001000100000: out_v[9] = 10'b1111100110;
    16'b0000101001000000: out_v[9] = 10'b0000001010;
    16'b1000101000000000: out_v[9] = 10'b1001001100;
    16'b0000100001100000: out_v[9] = 10'b0110100000;
    16'b0000001000000000: out_v[9] = 10'b0110111001;
    16'b1000100000000000: out_v[9] = 10'b1001001111;
    16'b1000001001000000: out_v[9] = 10'b0111111010;
    16'b1000000001000000: out_v[9] = 10'b1110010010;
    16'b0001001000000000: out_v[9] = 10'b0000101100;
    16'b0001101000000000: out_v[9] = 10'b0010001011;
    16'b0000000000100000: out_v[9] = 10'b0010011010;
    16'b0000001001000000: out_v[9] = 10'b1101010100;
    16'b0000000001000000: out_v[9] = 10'b0001011100;
    16'b0000100001000000: out_v[9] = 10'b0011101011;
    16'b0001101001000000: out_v[9] = 10'b1010011010;
    16'b0000000001100000: out_v[9] = 10'b0101111000;
    16'b1000000001100000: out_v[9] = 10'b1000100100;
    16'b0000100010100000: out_v[9] = 10'b1010010000;
    16'b0000110010100000: out_v[9] = 10'b0011110010;
    16'b0000000010100000: out_v[9] = 10'b0101111000;
    16'b1100000000000000: out_v[9] = 10'b1110100111;
    16'b1000100100101000: out_v[9] = 10'b1111110000;
    16'b1000101100100000: out_v[9] = 10'b1011010110;
    16'b1000100000101000: out_v[9] = 10'b0111001011;
    16'b1000100000001000: out_v[9] = 10'b0111011010;
    16'b0001000100000000: out_v[9] = 10'b0100001110;
    16'b0000001001100000: out_v[9] = 10'b1011000111;
    default: out_v[9] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000000100000: out_v[10] = 10'b1010000001;
    16'b0001001000000000: out_v[10] = 10'b1001110100;
    16'b0001001100010000: out_v[10] = 10'b0000000111;
    16'b0001001100110000: out_v[10] = 10'b1110011001;
    16'b0000000000110000: out_v[10] = 10'b0100100100;
    16'b0001001100000000: out_v[10] = 10'b1001000001;
    16'b0001001100100000: out_v[10] = 10'b1001110111;
    16'b0000001000110000: out_v[10] = 10'b1000101011;
    16'b0001000000100000: out_v[10] = 10'b0110001011;
    16'b0001001000100000: out_v[10] = 10'b0101100010;
    16'b0001000000000000: out_v[10] = 10'b1110001110;
    16'b0000001100100000: out_v[10] = 10'b1100010110;
    16'b0001001000110000: out_v[10] = 10'b0111101001;
    16'b0001001100100010: out_v[10] = 10'b0011001101;
    16'b0000001000010000: out_v[10] = 10'b0100110101;
    16'b0000001100110000: out_v[10] = 10'b1100000001;
    16'b0000001000100000: out_v[10] = 10'b0111011001;
    16'b0001001100000010: out_v[10] = 10'b1100000001;
    16'b1001000000100000: out_v[10] = 10'b0000000111;
    16'b0000000000000000: out_v[10] = 10'b1001010111;
    16'b0000001100000000: out_v[10] = 10'b0000110001;
    16'b0000001000000000: out_v[10] = 10'b0110110000;
    16'b1001000000000000: out_v[10] = 10'b1011001001;
    16'b0001001000010000: out_v[10] = 10'b0011111011;
    16'b0001000000110000: out_v[10] = 10'b0000100111;
    16'b0000001100010000: out_v[10] = 10'b0010011000;
    16'b0001000000000010: out_v[10] = 10'b1011110100;
    16'b1000000000000000: out_v[10] = 10'b0100111010;
    16'b1000000000000010: out_v[10] = 10'b1111110010;
    16'b1000000000100000: out_v[10] = 10'b0110010010;
    16'b1001001100100000: out_v[10] = 10'b1110000111;
    16'b1001000000110000: out_v[10] = 10'b0100101101;
    16'b1001000000010000: out_v[10] = 10'b0110000111;
    16'b1000001100000000: out_v[10] = 10'b0111100110;
    16'b1000000000110000: out_v[10] = 10'b0110000110;
    16'b0001000000110010: out_v[10] = 10'b0111110110;
    16'b0001000000010000: out_v[10] = 10'b1011010000;
    16'b0001000100110000: out_v[10] = 10'b0001101101;
    16'b1000001100100000: out_v[10] = 10'b0101100110;
    16'b1000000100100000: out_v[10] = 10'b1101101011;
    16'b0001000100100000: out_v[10] = 10'b0010001010;
    16'b0000000000010000: out_v[10] = 10'b0000110110;
    16'b1000000000010000: out_v[10] = 10'b0000111011;
    16'b1001000100110000: out_v[10] = 10'b0011111010;
    16'b0000000100000000: out_v[10] = 10'b0001100101;
    16'b1001000100100000: out_v[10] = 10'b1010101001;
    16'b1001000100000000: out_v[10] = 10'b0110101100;
    16'b1000000100000000: out_v[10] = 10'b0011100100;
    16'b1001000000100010: out_v[10] = 10'b0000111110;
    16'b0000000100100000: out_v[10] = 10'b0011011011;
    16'b1001001000100000: out_v[10] = 10'b0011111110;
    16'b1001001100110000: out_v[10] = 10'b0001010111;
    16'b0001000100000000: out_v[10] = 10'b0010101010;
    16'b0001000000100010: out_v[10] = 10'b0110011010;
    16'b0000000000110010: out_v[10] = 10'b1000111111;
    16'b1001000000110010: out_v[10] = 10'b1000010101;
    16'b1000000000110010: out_v[10] = 10'b0001001001;
    16'b1001000000000010: out_v[10] = 10'b0100011111;
    16'b0000000000100010: out_v[10] = 10'b1111100000;
    16'b1000001000110000: out_v[10] = 10'b1110000001;
    16'b1000001000010000: out_v[10] = 10'b1000110001;
    16'b1001001100000000: out_v[10] = 10'b0101010001;
    16'b1001001000000000: out_v[10] = 10'b1101100000;
    16'b1001001000010000: out_v[10] = 10'b0100110110;
    16'b1000001000000000: out_v[10] = 10'b0000011110;
    16'b1000001100010000: out_v[10] = 10'b1011010110;
    16'b1001001100010000: out_v[10] = 10'b1011001000;
    16'b1001001000110000: out_v[10] = 10'b1111000000;
    16'b0011001000010000: out_v[10] = 10'b1110000111;
    16'b0011000000010000: out_v[10] = 10'b1101101010;
    16'b1011001000010000: out_v[10] = 10'b0111111011;
    16'b0001000010010000: out_v[10] = 10'b1000010001;
    16'b0001000010000000: out_v[10] = 10'b0001001010;
    16'b0001001010000000: out_v[10] = 10'b1111010100;
    16'b0001001010010000: out_v[10] = 10'b0011111111;
    16'b0000000000000010: out_v[10] = 10'b1111101000;
    16'b1001000010000000: out_v[10] = 10'b1001101101;
    16'b1001001010000000: out_v[10] = 10'b1100010110;
    default: out_v[10] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010010001010000: out_v[11] = 10'b1000011111;
    16'b0010010100010100: out_v[11] = 10'b1100110101;
    16'b0011010100010100: out_v[11] = 10'b1011110111;
    16'b0011000011010100: out_v[11] = 10'b1110101011;
    16'b0010000011010000: out_v[11] = 10'b0010110011;
    16'b0010010000010000: out_v[11] = 10'b1101000000;
    16'b0011000000010000: out_v[11] = 10'b1001100100;
    16'b0010010100010000: out_v[11] = 10'b1111010100;
    16'b0011000111010100: out_v[11] = 10'b0001101010;
    16'b0010010011010000: out_v[11] = 10'b1010101110;
    16'b0010010010010100: out_v[11] = 10'b1110110100;
    16'b0010010110010100: out_v[11] = 10'b0011110110;
    16'b0011010101010100: out_v[11] = 10'b1111100010;
    16'b0010000001000100: out_v[11] = 10'b1101010001;
    16'b0011000001010100: out_v[11] = 10'b0010011010;
    16'b0010000111010100: out_v[11] = 10'b1001110111;
    16'b0010010001010100: out_v[11] = 10'b0101100100;
    16'b0010000011010100: out_v[11] = 10'b0110110011;
    16'b0010010011010100: out_v[11] = 10'b0111011100;
    16'b0011000011010000: out_v[11] = 10'b0001100011;
    16'b0010000101010100: out_v[11] = 10'b1011000111;
    16'b0001000001010000: out_v[11] = 10'b0001011011;
    16'b0011000101010100: out_v[11] = 10'b0110111010;
    16'b0001000001000100: out_v[11] = 10'b0011001001;
    16'b0011010011010100: out_v[11] = 10'b0011000100;
    16'b0000010000010100: out_v[11] = 10'b1010100011;
    16'b0000010010010100: out_v[11] = 10'b0010100011;
    16'b0010000010010100: out_v[11] = 10'b1001011011;
    16'b0011000001010000: out_v[11] = 10'b0010111001;
    16'b0010000100010100: out_v[11] = 10'b0111110011;
    16'b0001000011010000: out_v[11] = 10'b1110000011;
    16'b0011000101010000: out_v[11] = 10'b1111000001;
    16'b0010010000010100: out_v[11] = 10'b1110110010;
    16'b0011000001000100: out_v[11] = 10'b1101001101;
    16'b0010000100010000: out_v[11] = 10'b0111000011;
    16'b0010000001010100: out_v[11] = 10'b0110011011;
    16'b0011010001010100: out_v[11] = 10'b1111110010;
    16'b0010000001010000: out_v[11] = 10'b1001011011;
    16'b0010010111010100: out_v[11] = 10'b1111101100;
    16'b0010010010010000: out_v[11] = 10'b1001011100;
    16'b0011000101000100: out_v[11] = 10'b1001010111;
    16'b0000010100010000: out_v[11] = 10'b0000110111;
    16'b0010010101010100: out_v[11] = 10'b1111100000;
    16'b0010010000000100: out_v[11] = 10'b1010101111;
    16'b0001000001010100: out_v[11] = 10'b1011111101;
    16'b0011010111010100: out_v[11] = 10'b1100011101;
    16'b0011010001010000: out_v[11] = 10'b1010011110;
    16'b0001000011010100: out_v[11] = 10'b1111011010;
    16'b0000001000011101: out_v[11] = 10'b0110000110;
    16'b0000000000001000: out_v[11] = 10'b0111101011;
    16'b0000001000011001: out_v[11] = 10'b0100010011;
    16'b0000001010011001: out_v[11] = 10'b1110110000;
    16'b0000001000011000: out_v[11] = 10'b1010100110;
    16'b0000011001001000: out_v[11] = 10'b0001010011;
    16'b0000001000001101: out_v[11] = 10'b1111100011;
    16'b0000010001001000: out_v[11] = 10'b1000011101;
    16'b0000011000011001: out_v[11] = 10'b1100011110;
    16'b0000011010011001: out_v[11] = 10'b1011001001;
    16'b0000000001001000: out_v[11] = 10'b1011100001;
    16'b0000000001011000: out_v[11] = 10'b0011001001;
    16'b0000011001001001: out_v[11] = 10'b0010010011;
    16'b0000001010011000: out_v[11] = 10'b0110111000;
    16'b0000011001011000: out_v[11] = 10'b0100011011;
    16'b0000011000011101: out_v[11] = 10'b0000111110;
    16'b0000001010011101: out_v[11] = 10'b0010110011;
    16'b0000011000001101: out_v[11] = 10'b0010110000;
    16'b0000000010011000: out_v[11] = 10'b0110001110;
    16'b0000001000001001: out_v[11] = 10'b0001111101;
    16'b0000011010011101: out_v[11] = 10'b1010000010;
    16'b0000000000011000: out_v[11] = 10'b0011100011;
    16'b0000010000001000: out_v[11] = 10'b0010111101;
    16'b0000011000011000: out_v[11] = 10'b0001011001;
    16'b0000000010001000: out_v[11] = 10'b1011001101;
    16'b0000011011011001: out_v[11] = 10'b1111000011;
    16'b0000011000001000: out_v[11] = 10'b1000110000;
    16'b0000011001011001: out_v[11] = 10'b0110110010;
    16'b0000001001011001: out_v[11] = 10'b1010100100;
    16'b0011001001011001: out_v[11] = 10'b0100110110;
    16'b0000001011011101: out_v[11] = 10'b1001100100;
    16'b0010001000001001: out_v[11] = 10'b1011101011;
    16'b0001001011011101: out_v[11] = 10'b0111110100;
    16'b0010001011001001: out_v[11] = 10'b0111000101;
    16'b0010001011011001: out_v[11] = 10'b0101010100;
    16'b0011001011011001: out_v[11] = 10'b1111000100;
    16'b0010001010011001: out_v[11] = 10'b1110110010;
    16'b0010001011011000: out_v[11] = 10'b0011111011;
    16'b0011001001011000: out_v[11] = 10'b1010001110;
    16'b0000001011011001: out_v[11] = 10'b0101110101;
    16'b0011001010011000: out_v[11] = 10'b0111011111;
    16'b0011001010001001: out_v[11] = 10'b0111011100;
    16'b0011001011001001: out_v[11] = 10'b1100110010;
    16'b0011001011011101: out_v[11] = 10'b1011010110;
    16'b0011001010011001: out_v[11] = 10'b0111001001;
    16'b0010001001001001: out_v[11] = 10'b1010001101;
    16'b0000000001011100: out_v[11] = 10'b0111110001;
    16'b0011001000001001: out_v[11] = 10'b0001011101;
    16'b0011001001001001: out_v[11] = 10'b1000001000;
    16'b0000001011011000: out_v[11] = 10'b1010101111;
    16'b0000000011011100: out_v[11] = 10'b0100110110;
    16'b0010001010001001: out_v[11] = 10'b0111111111;
    16'b0000001011001001: out_v[11] = 10'b0001101111;
    16'b0011001011011000: out_v[11] = 10'b1011111001;
    16'b0000001011011100: out_v[11] = 10'b0011111111;
    16'b0001001001011001: out_v[11] = 10'b0110010111;
    16'b0010001001011001: out_v[11] = 10'b0110011101;
    16'b0000001001001001: out_v[11] = 10'b1001101101;
    16'b0011001001011101: out_v[11] = 10'b1010110111;
    16'b0000001010001001: out_v[11] = 10'b0010010000;
    16'b0011001011011100: out_v[11] = 10'b1010010110;
    16'b0001001011011001: out_v[11] = 10'b0011101000;
    16'b0000001001011101: out_v[11] = 10'b1010110101;
    16'b0010001011011101: out_v[11] = 10'b1000110111;
    16'b0010001011011100: out_v[11] = 10'b0010110100;
    16'b0011011001001001: out_v[11] = 10'b1110110101;
    16'b0010010001000100: out_v[11] = 10'b0100101010;
    16'b0011010001000100: out_v[11] = 10'b0010100010;
    16'b0010010001001100: out_v[11] = 10'b1011011111;
    16'b0010010001000000: out_v[11] = 10'b1000011101;
    16'b0010001001001100: out_v[11] = 10'b1110010010;
    16'b0000011001011100: out_v[11] = 10'b1001001111;
    16'b0010011001001100: out_v[11] = 10'b1111100101;
    16'b0001010001010000: out_v[11] = 10'b1010101010;
    16'b0000010001010000: out_v[11] = 10'b1000011100;
    16'b0000010011010100: out_v[11] = 10'b1001011110;
    16'b0010010001011100: out_v[11] = 10'b1010000111;
    16'b0001010001010100: out_v[11] = 10'b1010110110;
    16'b0010011001011100: out_v[11] = 10'b0001001111;
    16'b0011010011010000: out_v[11] = 10'b1010011000;
    16'b0000010011011100: out_v[11] = 10'b1011001100;
    16'b0011011001011000: out_v[11] = 10'b1001111000;
    16'b0001010001000100: out_v[11] = 10'b0101100111;
    16'b0000010001000100: out_v[11] = 10'b0101110010;
    16'b0000010001011100: out_v[11] = 10'b1000001101;
    16'b0000001001011100: out_v[11] = 10'b0000101111;
    16'b0000010001010100: out_v[11] = 10'b0101111011;
    16'b0011010001000000: out_v[11] = 10'b0000011110;
    16'b0010001001011100: out_v[11] = 10'b0011111111;
    16'b0010010011000100: out_v[11] = 10'b0001101101;
    16'b0010011011011100: out_v[11] = 10'b1011011011;
    16'b0010011001010100: out_v[11] = 10'b0010101110;
    16'b0011011001011100: out_v[11] = 10'b1011001101;
    16'b0010011001011000: out_v[11] = 10'b1011111010;
    16'b0000010001011000: out_v[11] = 10'b0101000101;
    16'b0000001000001000: out_v[11] = 10'b0001110111;
    16'b0000000001000000: out_v[11] = 10'b0110010101;
    16'b0000000000000000: out_v[11] = 10'b0111001010;
    16'b0000001001001000: out_v[11] = 10'b1010000101;
    16'b0010000000000000: out_v[11] = 10'b0110010000;
    16'b0000001001011000: out_v[11] = 10'b1011000001;
    16'b0000010000011000: out_v[11] = 10'b1001101010;
    16'b0011001000001000: out_v[11] = 10'b0001110111;
    16'b0000010000000000: out_v[11] = 10'b1101000110;
    16'b0010001000001000: out_v[11] = 10'b1000010011;
    16'b0000010000011100: out_v[11] = 10'b1001110101;
    16'b0010001001001000: out_v[11] = 10'b1001000001;
    16'b0000001000000000: out_v[11] = 10'b1101100010;
    16'b0000011000001001: out_v[11] = 10'b1000100100;
    16'b0010011001001001: out_v[11] = 10'b1010111100;
    16'b0010011000001000: out_v[11] = 10'b0001110010;
    16'b0000011000011100: out_v[11] = 10'b1010000101;
    16'b0000010001000000: out_v[11] = 10'b1110100100;
    16'b0010010000000000: out_v[11] = 10'b0000001101;
    16'b0010011000001001: out_v[11] = 10'b0111001100;
    16'b0000010100011000: out_v[11] = 10'b1001010101;
    16'b0000011100011000: out_v[11] = 10'b0110000010;
    16'b0000010000010000: out_v[11] = 10'b0010110100;
    16'b0000010100011100: out_v[11] = 10'b0111111110;
    16'b0000010100001000: out_v[11] = 10'b1000101010;
    16'b0000011100011100: out_v[11] = 10'b1001110001;
    16'b0000010100010100: out_v[11] = 10'b1010110111;
    16'b0000010100000000: out_v[11] = 10'b0001101011;
    16'b0001010011010000: out_v[11] = 10'b1101100110;
    16'b0010011011010001: out_v[11] = 10'b1101000010;
    16'b0010010010011000: out_v[11] = 10'b1111000110;
    16'b0010011011011001: out_v[11] = 10'b1111010010;
    16'b0000011010010000: out_v[11] = 10'b0110000111;
    16'b0010010011011000: out_v[11] = 10'b1100101101;
    16'b0011011010011001: out_v[11] = 10'b1110111011;
    16'b0010010000011000: out_v[11] = 10'b0111000111;
    16'b0010011010011000: out_v[11] = 10'b1001001011;
    16'b0010011001011001: out_v[11] = 10'b0101000010;
    16'b0010011010011001: out_v[11] = 10'b1010110011;
    16'b0011011011011001: out_v[11] = 10'b1110000001;
    16'b0010011000011001: out_v[11] = 10'b0111011010;
    16'b0010000001011000: out_v[11] = 10'b1111000101;
    16'b0010011011010000: out_v[11] = 10'b1011001100;
    16'b0011000011011000: out_v[11] = 10'b1111011010;
    16'b0010011011011000: out_v[11] = 10'b0010101010;
    16'b0000011010010001: out_v[11] = 10'b0011110101;
    16'b0000010010011000: out_v[11] = 10'b1101001100;
    16'b0010011000011000: out_v[11] = 10'b1100100000;
    16'b0010011010010000: out_v[11] = 10'b1011001110;
    16'b0010000011011000: out_v[11] = 10'b0101010111;
    16'b0010011010010001: out_v[11] = 10'b1011011100;
    16'b0010000000011000: out_v[11] = 10'b1101001000;
    16'b0010011010001001: out_v[11] = 10'b0011101011;
    16'b0010000001001000: out_v[11] = 10'b0111001010;
    16'b0011000000011000: out_v[11] = 10'b1110101011;
    16'b0011000001011000: out_v[11] = 10'b1100101100;
    16'b0011011001011001: out_v[11] = 10'b1101011100;
    16'b0000011010011000: out_v[11] = 10'b1110101101;
    16'b0000000000010000: out_v[11] = 10'b1000101110;
    16'b0010000000010000: out_v[11] = 10'b0110111010;
    16'b0000000000011100: out_v[11] = 10'b0010100010;
    16'b0000000001010000: out_v[11] = 10'b1110110110;
    16'b0000000000010100: out_v[11] = 10'b1111010001;
    16'b0000000100011100: out_v[11] = 10'b0011001000;
    16'b0000000100010100: out_v[11] = 10'b1011101110;
    16'b0000011001001100: out_v[11] = 10'b1111000110;
    16'b0000011001001101: out_v[11] = 10'b1001010011;
    16'b0000011001011101: out_v[11] = 10'b1101011000;
    16'b0000011011011101: out_v[11] = 10'b1110001000;
    16'b0000001100011101: out_v[11] = 10'b1111001000;
    16'b0000001001001101: out_v[11] = 10'b0111010011;
    16'b0000011101001101: out_v[11] = 10'b1010101111;
    16'b0000011101011101: out_v[11] = 10'b1001111100;
    16'b0010011001011101: out_v[11] = 10'b1111100101;
    16'b0000011100011101: out_v[11] = 10'b0011111100;
    16'b0000011100001101: out_v[11] = 10'b1011010010;
    16'b0000011101011100: out_v[11] = 10'b0001100111;
    16'b0010011011011101: out_v[11] = 10'b1001001100;
    16'b0010011001001101: out_v[11] = 10'b0011100011;
    16'b0000001101011101: out_v[11] = 10'b1001110110;
    16'b0000001101001101: out_v[11] = 10'b0111110011;
    16'b0010011001010001: out_v[11] = 10'b0100110001;
    16'b0000001000010000: out_v[11] = 10'b0111111101;
    16'b0000001000011100: out_v[11] = 10'b0101111001;
    16'b0010000001000000: out_v[11] = 10'b0010100010;
    16'b0000001001000000: out_v[11] = 10'b1000110111;
    16'b0010001000000000: out_v[11] = 10'b1001011011;
    16'b0000011000000000: out_v[11] = 10'b1010000111;
    default: out_v[11] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000000001000: out_v[12] = 10'b0000110110;
    16'b0000000011000000: out_v[12] = 10'b0100011100;
    16'b0010000001001000: out_v[12] = 10'b0001001001;
    16'b1000000001001000: out_v[12] = 10'b0011001001;
    16'b1000000011001000: out_v[12] = 10'b1001000100;
    16'b0110000001001000: out_v[12] = 10'b1101100011;
    16'b0000000011001000: out_v[12] = 10'b1001000101;
    16'b1000000001000000: out_v[12] = 10'b0101000011;
    16'b0000000001001000: out_v[12] = 10'b1001011111;
    16'b0000000010001000: out_v[12] = 10'b0000011110;
    16'b0000000000000000: out_v[12] = 10'b1001110111;
    16'b0100000001001000: out_v[12] = 10'b0100101011;
    16'b0000000001000000: out_v[12] = 10'b1000001111;
    16'b1000000010001000: out_v[12] = 10'b0100010101;
    16'b1000000011000000: out_v[12] = 10'b0111001110;
    16'b0010000011001000: out_v[12] = 10'b0011011110;
    16'b0110000011001000: out_v[12] = 10'b1001001010;
    16'b1110000001001000: out_v[12] = 10'b1110100011;
    16'b0000000010000000: out_v[12] = 10'b1001010100;
    16'b0110000001000000: out_v[12] = 10'b1100110000;
    16'b0110000000001000: out_v[12] = 10'b1001101011;
    16'b0010000001000000: out_v[12] = 10'b0011100010;
    16'b0100000011001000: out_v[12] = 10'b1011101110;
    16'b1010000001001000: out_v[12] = 10'b0010110110;
    16'b1000000000001000: out_v[12] = 10'b1000110110;
    16'b1000000010000000: out_v[12] = 10'b0111100100;
    16'b1000000000000000: out_v[12] = 10'b0100111010;
    16'b0010000000001000: out_v[12] = 10'b1000001110;
    16'b0010000000000000: out_v[12] = 10'b0100001110;
    16'b0010000010000000: out_v[12] = 10'b1110000000;
    16'b0010000010001000: out_v[12] = 10'b0100000110;
    16'b1010000000001000: out_v[12] = 10'b0010100111;
    16'b0010000011000000: out_v[12] = 10'b0011010011;
    16'b0110000011000000: out_v[12] = 10'b1100010001;
    16'b0100000011000000: out_v[12] = 10'b0011110011;
    16'b0100000001000000: out_v[12] = 10'b0011111010;
    16'b0010000010010010: out_v[12] = 10'b0101010011;
    16'b0110000000000000: out_v[12] = 10'b1111001001;
    16'b0000000010010010: out_v[12] = 10'b1100000010;
    16'b0010000000010010: out_v[12] = 10'b0111110011;
    16'b0000000000010000: out_v[12] = 10'b0010101111;
    16'b0000000001010010: out_v[12] = 10'b1001101110;
    16'b0000000000010010: out_v[12] = 10'b1011101101;
    16'b0100000000000000: out_v[12] = 10'b1110001110;
    16'b0110000010000000: out_v[12] = 10'b1010011101;
    16'b0000000011010010: out_v[12] = 10'b0111000111;
    16'b0110000010010010: out_v[12] = 10'b0011111000;
    16'b0100000010000000: out_v[12] = 10'b0011100110;
    default: out_v[12] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000100000100: out_v[13] = 10'b0001110001;
    16'b0000000100110110: out_v[13] = 10'b0010001001;
    16'b0000000100110100: out_v[13] = 10'b1010110010;
    16'b0000000000110110: out_v[13] = 10'b1110010001;
    16'b0000000000110010: out_v[13] = 10'b0011000000;
    16'b0000000000110000: out_v[13] = 10'b0000011001;
    16'b0000000100010011: out_v[13] = 10'b0011111001;
    16'b0000000100110000: out_v[13] = 10'b1000011011;
    16'b0000000100010110: out_v[13] = 10'b0010010101;
    16'b0000000100110111: out_v[13] = 10'b0101100101;
    16'b0000000000110100: out_v[13] = 10'b1010010001;
    16'b0000000100010111: out_v[13] = 10'b0011010111;
    16'b0000000100000110: out_v[13] = 10'b1000110101;
    16'b0000100000110110: out_v[13] = 10'b0100011111;
    16'b0000000100110010: out_v[13] = 10'b1001011000;
    16'b0000000100000010: out_v[13] = 10'b0001101111;
    16'b0000100100110110: out_v[13] = 10'b1001111010;
    16'b0000000100100100: out_v[13] = 10'b0011000011;
    16'b0000000100000111: out_v[13] = 10'b0101010001;
    16'b0000000100010100: out_v[13] = 10'b0000111111;
    16'b0000100000110100: out_v[13] = 10'b0011110110;
    16'b0000000000010010: out_v[13] = 10'b1011011000;
    16'b0000000100010010: out_v[13] = 10'b0110110001;
    16'b0000000000010110: out_v[13] = 10'b0101011111;
    16'b0001100000000000: out_v[13] = 10'b1011111010;
    16'b0001100000010000: out_v[13] = 10'b0010110010;
    16'b0001000100010000: out_v[13] = 10'b0100010010;
    16'b0001000000010000: out_v[13] = 10'b1011000001;
    16'b0001000100110000: out_v[13] = 10'b1010100011;
    16'b0001000100100000: out_v[13] = 10'b1110100000;
    16'b0001100100010000: out_v[13] = 10'b0101010110;
    16'b0001100000110000: out_v[13] = 10'b0101000001;
    16'b0001000000000000: out_v[13] = 10'b1000001111;
    16'b0001000100000000: out_v[13] = 10'b0101111000;
    16'b0001100000000100: out_v[13] = 10'b1010111010;
    16'b0001000000100000: out_v[13] = 10'b1011000111;
    16'b0001000000110000: out_v[13] = 10'b1000101111;
    16'b0001100100110000: out_v[13] = 10'b0111010000;
    16'b0001100100010001: out_v[13] = 10'b1101000101;
    16'b0001100000110001: out_v[13] = 10'b0000000101;
    16'b0001000000110101: out_v[13] = 10'b1011101111;
    16'b0001000000000100: out_v[13] = 10'b1110001011;
    16'b0001100000100000: out_v[13] = 10'b0001001101;
    16'b0001000100010001: out_v[13] = 10'b1010011001;
    16'b0001000000110001: out_v[13] = 10'b1101111010;
    16'b0001100000000110: out_v[13] = 10'b1011010110;
    16'b0001100000110100: out_v[13] = 10'b1111001000;
    16'b0001100000100110: out_v[13] = 10'b0001100110;
    16'b0000100000110000: out_v[13] = 10'b0001110010;
    16'b0001100000100100: out_v[13] = 10'b0011100101;
    16'b0001000000110111: out_v[13] = 10'b1001000100;
    16'b0001100000100001: out_v[13] = 10'b0001101101;
    16'b0000100000110001: out_v[13] = 10'b0111001011;
    16'b0001000000010001: out_v[13] = 10'b0010100101;
    16'b0001100000000001: out_v[13] = 10'b1010011110;
    16'b0000000000110001: out_v[13] = 10'b1110011010;
    16'b0001000000110100: out_v[13] = 10'b1101001100;
    16'b0000100000100100: out_v[13] = 10'b1001111000;
    16'b0000100000110101: out_v[13] = 10'b0001101100;
    16'b0000100000100000: out_v[13] = 10'b0010111000;
    16'b0001100000110101: out_v[13] = 10'b1011111011;
    16'b0001100000010001: out_v[13] = 10'b1110000101;
    16'b0001100100010101: out_v[13] = 10'b1001010111;
    16'b0001100100010100: out_v[13] = 10'b0111100100;
    16'b0001000000110110: out_v[13] = 10'b0101000110;
    16'b0001100100110001: out_v[13] = 10'b1100010101;
    16'b0001100000100101: out_v[13] = 10'b0101001111;
    16'b0001000000100100: out_v[13] = 10'b0111110010;
    16'b0001100000010100: out_v[13] = 10'b0111111011;
    16'b0000000100000000: out_v[13] = 10'b0101100101;
    16'b0001000100110001: out_v[13] = 10'b0010100100;
    16'b0001000100001001: out_v[13] = 10'b1111001111;
    16'b0001000100100100: out_v[13] = 10'b0100010001;
    16'b0000000100010001: out_v[13] = 10'b1100010110;
    16'b0001000100000101: out_v[13] = 10'b0101001011;
    16'b0000000100000001: out_v[13] = 10'b1101110111;
    16'b0000000100100000: out_v[13] = 10'b1011100011;
    16'b0001000100000001: out_v[13] = 10'b1011100011;
    16'b0001000100110100: out_v[13] = 10'b0010101010;
    16'b0001000100110101: out_v[13] = 10'b1101011011;
    16'b0000000100110001: out_v[13] = 10'b0111010100;
    16'b0000000100100001: out_v[13] = 10'b0111110110;
    16'b0000000100010000: out_v[13] = 10'b1001010100;
    16'b0001000100010011: out_v[13] = 10'b0000111010;
    16'b0001000100000100: out_v[13] = 10'b0110001110;
    16'b0001000100100001: out_v[13] = 10'b1000101001;
    16'b0001000100010101: out_v[13] = 10'b0010001100;
    16'b0000000100110101: out_v[13] = 10'b1100010100;
    16'b0001000100010100: out_v[13] = 10'b0011011010;
    16'b0001000000010010: out_v[13] = 10'b0101011000;
    16'b0001000000100010: out_v[13] = 10'b0011011010;
    16'b0001100000010010: out_v[13] = 10'b0101010001;
    16'b0001000000100111: out_v[13] = 10'b1011111001;
    16'b0001100000010110: out_v[13] = 10'b0010011010;
    16'b0001000100100110: out_v[13] = 10'b1100000000;
    16'b0001000100100010: out_v[13] = 10'b0111010011;
    16'b0001000000010110: out_v[13] = 10'b1101100001;
    16'b0001000000000110: out_v[13] = 10'b1001110001;
    16'b0001000000000111: out_v[13] = 10'b0000010010;
    16'b0000000100100110: out_v[13] = 10'b0011001110;
    16'b0001000100100111: out_v[13] = 10'b1110000111;
    16'b0001000000100011: out_v[13] = 10'b0110000101;
    16'b0001000000100110: out_v[13] = 10'b1001110110;
    16'b0001000000000010: out_v[13] = 10'b1010100110;
    16'b0001000000010100: out_v[13] = 10'b0100010001;
    16'b0001000100110110: out_v[13] = 10'b1001110111;
    16'b0000100100100000: out_v[13] = 10'b1000111010;
    16'b0001000000110010: out_v[13] = 10'b0001001100;
    16'b0001100000110110: out_v[13] = 10'b0011011001;
    16'b0001100000000010: out_v[13] = 10'b1100001000;
    16'b0001000000000011: out_v[13] = 10'b1111001010;
    16'b0001000100110010: out_v[13] = 10'b0010101101;
    16'b0001000100100011: out_v[13] = 10'b1101011011;
    16'b0000100000100110: out_v[13] = 10'b0100011011;
    16'b0000000000010000: out_v[13] = 10'b1110100001;
    16'b0001000100000010: out_v[13] = 10'b0111110110;
    16'b0000000000000000: out_v[13] = 10'b0010110010;
    16'b0000100000010000: out_v[13] = 10'b1100101000;
    16'b0001000100010010: out_v[13] = 10'b1001101110;
    16'b0001100000110010: out_v[13] = 10'b0111011011;
    16'b0001100000110011: out_v[13] = 10'b1111001111;
    16'b0001100000110111: out_v[13] = 10'b1001010110;
    16'b0000100000110010: out_v[13] = 10'b1111000100;
    16'b0001100000100010: out_v[13] = 10'b1101001101;
    16'b0001100000100111: out_v[13] = 10'b1110111011;
    16'b0000000000100000: out_v[13] = 10'b0011110111;
    16'b0000000000000110: out_v[13] = 10'b0010010010;
    16'b0000000000010100: out_v[13] = 10'b1110000001;
    16'b0000000000000100: out_v[13] = 10'b1010100110;
    16'b0000000100100010: out_v[13] = 10'b1111001110;
    16'b0001100100110101: out_v[13] = 10'b0101001000;
    16'b0001100100100100: out_v[13] = 10'b0111001011;
    16'b0001100100110100: out_v[13] = 10'b0100101110;
    16'b0001100100100000: out_v[13] = 10'b1110001001;
    16'b0001100100000100: out_v[13] = 10'b0100110111;
    16'b0001100100000000: out_v[13] = 10'b0111001101;
    16'b0001100100110110: out_v[13] = 10'b1101000010;
    16'b0000100100100110: out_v[13] = 10'b0101111101;
    16'b0001100100100110: out_v[13] = 10'b1100100011;
    16'b0000100000000110: out_v[13] = 10'b1100001011;
    default: out_v[13] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100000110000000: out_v[14] = 10'b0100100100;
    16'b0100000100000000: out_v[14] = 10'b1110000001;
    16'b0110001110000000: out_v[14] = 10'b1111010011;
    16'b0100000010000000: out_v[14] = 10'b0110110001;
    16'b0100001011000000: out_v[14] = 10'b0111011011;
    16'b0110000010000000: out_v[14] = 10'b1011010100;
    16'b0000000000000000: out_v[14] = 10'b0010100010;
    16'b0000000110000000: out_v[14] = 10'b0011100111;
    16'b0000001110000000: out_v[14] = 10'b0101011011;
    16'b0100000110000001: out_v[14] = 10'b0100100001;
    16'b0100100110000001: out_v[14] = 10'b1110001000;
    16'b0100000010000001: out_v[14] = 10'b1000010111;
    16'b0100001110000000: out_v[14] = 10'b0011100010;
    16'b0100000000000000: out_v[14] = 10'b1010010100;
    16'b0110000110000000: out_v[14] = 10'b0111101110;
    16'b0000000010000000: out_v[14] = 10'b1000110101;
    16'b0100001111000000: out_v[14] = 10'b1001101101;
    16'b0000000010000001: out_v[14] = 10'b0000101110;
    16'b0000001111000000: out_v[14] = 10'b0100010101;
    16'b0100001100000000: out_v[14] = 10'b0110110001;
    16'b0110001010000000: out_v[14] = 10'b0111101010;
    16'b0000000110000001: out_v[14] = 10'b0011101001;
    16'b0100001001000000: out_v[14] = 10'b0010011001;
    16'b0000000100000000: out_v[14] = 10'b0010110111;
    16'b0000001100000000: out_v[14] = 10'b0100110111;
    16'b0100000100000001: out_v[14] = 10'b1100110011;
    16'b0110000100000000: out_v[14] = 10'b0010011010;
    16'b0010000010000000: out_v[14] = 10'b1100010101;
    16'b0100100110000000: out_v[14] = 10'b0110110101;
    16'b0000001011000000: out_v[14] = 10'b1101011100;
    16'b0110000010000001: out_v[14] = 10'b0100101111;
    16'b0000000100000001: out_v[14] = 10'b0111011000;
    16'b0110000110000001: out_v[14] = 10'b1100011011;
    16'b0100001010000000: out_v[14] = 10'b0100011111;
    16'b0100001000000000: out_v[14] = 10'b1001110100;
    16'b0000100010000001: out_v[14] = 10'b0011110000;
    16'b0000100100000001: out_v[14] = 10'b1101001010;
    16'b0000100000000001: out_v[14] = 10'b1000100000;
    16'b0000000000000001: out_v[14] = 10'b1101001010;
    16'b0000100100000000: out_v[14] = 10'b0010010011;
    16'b0000100110000001: out_v[14] = 10'b0111000000;
    16'b0000100010000000: out_v[14] = 10'b0010110110;
    16'b0000100000000000: out_v[14] = 10'b0110010000;
    16'b0000100110000000: out_v[14] = 10'b1101000111;
    16'b0000101011000001: out_v[14] = 10'b1011100111;
    16'b0001100010000001: out_v[14] = 10'b0111111011;
    16'b0000101000000001: out_v[14] = 10'b1110101110;
    16'b0110100000000001: out_v[14] = 10'b0010001110;
    16'b0000101001000000: out_v[14] = 10'b0100111011;
    16'b0100100010000000: out_v[14] = 10'b1011001000;
    16'b0000101010000000: out_v[14] = 10'b1000000101;
    16'b0101000010000000: out_v[14] = 10'b1110111011;
    16'b0110000000000000: out_v[14] = 10'b1100010110;
    16'b0000101011000000: out_v[14] = 10'b1011000011;
    16'b0000001001000001: out_v[14] = 10'b1110110110;
    16'b0100100010000001: out_v[14] = 10'b1001010110;
    16'b0000101001000001: out_v[14] = 10'b0101111110;
    16'b0110100000000000: out_v[14] = 10'b1100110011;
    16'b0000101000000000: out_v[14] = 10'b1100010010;
    16'b0001100010000000: out_v[14] = 10'b0011001101;
    16'b0100100000000000: out_v[14] = 10'b1001100010;
    16'b0000101010000001: out_v[14] = 10'b1010001000;
    16'b0001100000000000: out_v[14] = 10'b0101001111;
    16'b0100100100000001: out_v[14] = 10'b0110010000;
    16'b0000101110000001: out_v[14] = 10'b1101011000;
    16'b0010100110000001: out_v[14] = 10'b1110110101;
    16'b0110100010000001: out_v[14] = 10'b0100011010;
    16'b0100101100000001: out_v[14] = 10'b1100001000;
    16'b0000101100000001: out_v[14] = 10'b0010001011;
    16'b0010100010000001: out_v[14] = 10'b0011000111;
    16'b0110100110000001: out_v[14] = 10'b1001101010;
    16'b0100101110000001: out_v[14] = 10'b0110011010;
    16'b0100000000000001: out_v[14] = 10'b1001001110;
    16'b0100100100000000: out_v[14] = 10'b1010111111;
    16'b0100100000000001: out_v[14] = 10'b0100011111;
    16'b0000001000000000: out_v[14] = 10'b1011101011;
    16'b0000000010100000: out_v[14] = 10'b1100110111;
    16'b0100100010100001: out_v[14] = 10'b0011110110;
    16'b0000000010100001: out_v[14] = 10'b1011001000;
    16'b0101100000000001: out_v[14] = 10'b1111001111;
    16'b0101101001000000: out_v[14] = 10'b0001111100;
    16'b0101100000000000: out_v[14] = 10'b1101100011;
    16'b0000000000100000: out_v[14] = 10'b0111101011;
    16'b0100101000000000: out_v[14] = 10'b1011011010;
    16'b0100101000000001: out_v[14] = 10'b0110111010;
    16'b0000000000100001: out_v[14] = 10'b1001110001;
    16'b0000100010100001: out_v[14] = 10'b0000110010;
    16'b0100101001000001: out_v[14] = 10'b0111101000;
    16'b0100000000000010: out_v[14] = 10'b0000010111;
    16'b0000100000000010: out_v[14] = 10'b0011100011;
    16'b0100000100000010: out_v[14] = 10'b0110000010;
    16'b0000000000000010: out_v[14] = 10'b1101110010;
    16'b0100100100000010: out_v[14] = 10'b1111110110;
    default: out_v[14] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1010000110000000: out_v[15] = 10'b0100011001;
    16'b1010000111000000: out_v[15] = 10'b0101100000;
    16'b1110100110000000: out_v[15] = 10'b1001011001;
    16'b1000000110000000: out_v[15] = 10'b1010011101;
    16'b1110100000000000: out_v[15] = 10'b0110010001;
    16'b1010000101000000: out_v[15] = 10'b0011100000;
    16'b1010000000000000: out_v[15] = 10'b1100100001;
    16'b0000000110000000: out_v[15] = 10'b1110000110;
    16'b1010000100000000: out_v[15] = 10'b1111100000;
    16'b0100100110000000: out_v[15] = 10'b0111000011;
    16'b0010000111000000: out_v[15] = 10'b0100110101;
    16'b0010000110000000: out_v[15] = 10'b0101000011;
    16'b0010000011000000: out_v[15] = 10'b1110001111;
    16'b1110100100000000: out_v[15] = 10'b1101100011;
    16'b1010100100000000: out_v[15] = 10'b1100100010;
    16'b0000000111000000: out_v[15] = 10'b1001010111;
    16'b1010100110000000: out_v[15] = 10'b0100001110;
    16'b1100100100000000: out_v[15] = 10'b1100010010;
    16'b1010000010000000: out_v[15] = 10'b0100111011;
    16'b1100100110000000: out_v[15] = 10'b0100011100;
    16'b1110100111000000: out_v[15] = 10'b1011100111;
    16'b1000000100000000: out_v[15] = 10'b1101010010;
    16'b1010100000000000: out_v[15] = 10'b0111100100;
    16'b1000000000000000: out_v[15] = 10'b0000111011;
    16'b0010000000000000: out_v[15] = 10'b1010011011;
    16'b1000000010000000: out_v[15] = 10'b1000011011;
    16'b1110000110000000: out_v[15] = 10'b0111001100;
    16'b1000100110000000: out_v[15] = 10'b0000011111;
    16'b0010000101000000: out_v[15] = 10'b1000101101;
    16'b0010000010000000: out_v[15] = 10'b0011111000;
    16'b0110100110000000: out_v[15] = 10'b0111100001;
    16'b1110000100000000: out_v[15] = 10'b0010110110;
    16'b0000000000000000: out_v[15] = 10'b1011100010;
    16'b0000000010000000: out_v[15] = 10'b0000110000;
    16'b0010100000000000: out_v[15] = 10'b1000011111;
    16'b1000000101000000: out_v[15] = 10'b0001110010;
    16'b0110100000000000: out_v[15] = 10'b0000001010;
    16'b1100000000000000: out_v[15] = 10'b1011011110;
    16'b1100100010000000: out_v[15] = 10'b0101011100;
    16'b1110100010000000: out_v[15] = 10'b1111011001;
    16'b1100000110000000: out_v[15] = 10'b1010100111;
    16'b1110000000000000: out_v[15] = 10'b0000100110;
    16'b0100100000000000: out_v[15] = 10'b1001100000;
    16'b1100000010000000: out_v[15] = 10'b0110100111;
    16'b0110000000000000: out_v[15] = 10'b1010000110;
    16'b1000100100000000: out_v[15] = 10'b1111010110;
    16'b1000100000000000: out_v[15] = 10'b0111001100;
    16'b0000100010000000: out_v[15] = 10'b0111110010;
    16'b0100000000000000: out_v[15] = 10'b1001100101;
    16'b1000100010000000: out_v[15] = 10'b0100010101;
    16'b0000100000000000: out_v[15] = 10'b0011011011;
    16'b0110100010000000: out_v[15] = 10'b0101100010;
    16'b1000000111000000: out_v[15] = 10'b1010001011;
    16'b1010100010000000: out_v[15] = 10'b1000000111;
    16'b1000100111000000: out_v[15] = 10'b0111000101;
    16'b1010100111000000: out_v[15] = 10'b1011101110;
    16'b1010000100010000: out_v[15] = 10'b1000101010;
    16'b0010000000010000: out_v[15] = 10'b0110011001;
    16'b1010000000010000: out_v[15] = 10'b1001100000;
    16'b0010100010000000: out_v[15] = 10'b0110100110;
    16'b1000000101010000: out_v[15] = 10'b0000110000;
    16'b0000000101000000: out_v[15] = 10'b0010111101;
    16'b1000000100010000: out_v[15] = 10'b0110110101;
    16'b0000000001000000: out_v[15] = 10'b0000011111;
    16'b0010000100000000: out_v[15] = 10'b1100100010;
    16'b0010000101010000: out_v[15] = 10'b1100000111;
    16'b1010000101010000: out_v[15] = 10'b1110110110;
    16'b0100100010000000: out_v[15] = 10'b1011100010;
    16'b0100010000000000: out_v[15] = 10'b0101101111;
    16'b0100110000000000: out_v[15] = 10'b1111000001;
    16'b1000010000000000: out_v[15] = 10'b1111010001;
    16'b0000010000000000: out_v[15] = 10'b0101100011;
    16'b0110000010000000: out_v[15] = 10'b1011110110;
    16'b1000000000010000: out_v[15] = 10'b0010100111;
    16'b0010000100010000: out_v[15] = 10'b1100100110;
    default: out_v[15] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100000000010001: out_v[16] = 10'b0110000011;
    16'b0100000000010100: out_v[16] = 10'b0111011001;
    16'b0100100000010100: out_v[16] = 10'b0000111111;
    16'b0100101000000111: out_v[16] = 10'b0111110011;
    16'b0100000000010011: out_v[16] = 10'b1100101101;
    16'b0000000000010011: out_v[16] = 10'b0010110101;
    16'b0000100000010000: out_v[16] = 10'b1001110001;
    16'b0100101000000110: out_v[16] = 10'b1101011110;
    16'b0000100000000100: out_v[16] = 10'b0111000110;
    16'b0000100000010100: out_v[16] = 10'b0100000001;
    16'b0000101000000100: out_v[16] = 10'b0011001011;
    16'b0100000000010101: out_v[16] = 10'b0100011010;
    16'b0100000000000100: out_v[16] = 10'b1001100110;
    16'b0100100000000001: out_v[16] = 10'b1111111101;
    16'b0000000000010001: out_v[16] = 10'b1001101011;
    16'b0100101000000001: out_v[16] = 10'b0000011111;
    16'b0100100000010001: out_v[16] = 10'b1101001010;
    16'b0000100000000000: out_v[16] = 10'b0100110111;
    16'b0100100000000100: out_v[16] = 10'b1011010011;
    16'b0100000000000001: out_v[16] = 10'b1110011000;
    16'b0101100000010001: out_v[16] = 10'b0111011011;
    16'b0100100000010111: out_v[16] = 10'b0001111011;
    16'b0100001000000100: out_v[16] = 10'b1011100111;
    16'b0100100000000110: out_v[16] = 10'b1110110011;
    16'b0100101000000101: out_v[16] = 10'b0001011111;
    16'b0100101000000100: out_v[16] = 10'b0110110101;
    16'b0001100000010001: out_v[16] = 10'b0001110011;
    16'b0100100000000011: out_v[16] = 10'b0110100111;
    16'b0100000000010010: out_v[16] = 10'b0101000010;
    16'b0100100000010101: out_v[16] = 10'b1100010011;
    16'b0100100000010110: out_v[16] = 10'b1110111100;
    16'b0100101000000000: out_v[16] = 10'b1001001001;
    16'b0100100000000101: out_v[16] = 10'b1010000110;
    16'b0100000000010111: out_v[16] = 10'b1110110010;
    16'b0000100000010001: out_v[16] = 10'b1100110111;
    16'b0100000000010000: out_v[16] = 10'b0111010010;
    16'b0100100000000000: out_v[16] = 10'b0000111001;
    16'b0100000000000011: out_v[16] = 10'b1111101101;
    16'b0101100000010100: out_v[16] = 10'b1010001101;
    16'b0100000000010110: out_v[16] = 10'b1010111111;
    16'b0100101000000011: out_v[16] = 10'b1000000101;
    16'b0100100000010011: out_v[16] = 10'b0011100111;
    16'b0100000000000000: out_v[16] = 10'b0010101011;
    16'b0101100000000100: out_v[16] = 10'b0011101100;
    16'b0000100000010101: out_v[16] = 10'b1000101011;
    16'b0000000000000000: out_v[16] = 10'b1111001010;
    16'b0000000000000010: out_v[16] = 10'b0001100111;
    16'b0100000000000010: out_v[16] = 10'b0010100001;
    16'b0000000000010000: out_v[16] = 10'b0000111110;
    16'b0000001000010000: out_v[16] = 10'b0100110110;
    16'b0000000000010010: out_v[16] = 10'b0001001100;
    16'b0001000100000000: out_v[16] = 10'b0101011001;
    16'b0000000000000001: out_v[16] = 10'b1111010011;
    16'b0001000000010001: out_v[16] = 10'b0000001101;
    16'b0001000000000000: out_v[16] = 10'b1010110101;
    16'b0000001000010011: out_v[16] = 10'b1000001101;
    16'b0101000000000001: out_v[16] = 10'b0010011100;
    16'b0101000000010000: out_v[16] = 10'b1111110110;
    16'b0000101000010011: out_v[16] = 10'b0010111011;
    16'b0000001000010010: out_v[16] = 10'b0010010101;
    16'b0000100000000011: out_v[16] = 10'b1111001111;
    16'b0101000000000000: out_v[16] = 10'b1010001011;
    16'b0001000000000001: out_v[16] = 10'b0110101101;
    16'b0101000000010001: out_v[16] = 10'b0011101010;
    16'b0000001000000011: out_v[16] = 10'b1011110101;
    16'b0000000000000011: out_v[16] = 10'b0100001110;
    16'b0000100000010011: out_v[16] = 10'b0011101010;
    16'b0000001000010001: out_v[16] = 10'b1100010111;
    16'b0000001000010101: out_v[16] = 10'b0011010100;
    16'b0000000001010000: out_v[16] = 10'b0101101110;
    16'b0001000000010000: out_v[16] = 10'b1010101010;
    16'b0000101000000011: out_v[16] = 10'b1001001100;
    16'b0101000100010001: out_v[16] = 10'b0111010100;
    16'b0000001000000001: out_v[16] = 10'b1100101000;
    16'b0101000000010011: out_v[16] = 10'b1011101110;
    16'b0001000000010010: out_v[16] = 10'b1011011010;
    16'b0000001000010111: out_v[16] = 10'b1101111010;
    16'b0101001000000000: out_v[16] = 10'b1010101111;
    16'b0100001000000011: out_v[16] = 10'b1001110110;
    16'b0101001000000001: out_v[16] = 10'b1010101010;
    16'b0100001000000001: out_v[16] = 10'b1011110000;
    16'b0100001000000000: out_v[16] = 10'b0010101010;
    16'b0100001000000010: out_v[16] = 10'b0001111101;
    16'b0101000100000000: out_v[16] = 10'b0011101010;
    16'b0101000100000001: out_v[16] = 10'b1001101111;
    16'b0000001000000000: out_v[16] = 10'b1011111000;
    16'b0100001000000101: out_v[16] = 10'b0001001010;
    16'b0101001000000011: out_v[16] = 10'b1011111001;
    16'b0100000000000101: out_v[16] = 10'b0111011100;
    16'b0001100000000001: out_v[16] = 10'b0111010110;
    16'b0000000100000001: out_v[16] = 10'b1000010101;
    16'b0000000100000000: out_v[16] = 10'b1110000011;
    16'b0001100100010001: out_v[16] = 10'b1010100110;
    16'b0000100100000001: out_v[16] = 10'b0101010010;
    16'b0000100000000001: out_v[16] = 10'b0110111000;
    16'b0001000100000001: out_v[16] = 10'b1100101000;
    16'b0000100000000101: out_v[16] = 10'b0011001010;
    16'b0001100100000001: out_v[16] = 10'b1010100110;
    16'b0000100100010001: out_v[16] = 10'b1101001000;
    16'b0000000000000100: out_v[16] = 10'b0001110111;
    16'b0100000100000000: out_v[16] = 10'b1000001110;
    16'b0000000000010100: out_v[16] = 10'b0001101011;
    16'b0000010000010010: out_v[16] = 10'b1010110011;
    16'b0001000001010001: out_v[16] = 10'b1110111101;
    16'b0000010000010000: out_v[16] = 10'b0111011000;
    16'b0000000001010001: out_v[16] = 10'b0100100111;
    16'b0000100000010010: out_v[16] = 10'b0001011100;
    16'b0000000001000001: out_v[16] = 10'b1111100001;
    16'b0000000000010101: out_v[16] = 10'b0111001001;
    16'b0101000000000101: out_v[16] = 10'b1110001111;
    16'b0000000000000101: out_v[16] = 10'b0000111100;
    16'b0100001000010101: out_v[16] = 10'b0100010111;
    16'b0101000000010101: out_v[16] = 10'b1111000010;
    16'b0100001000010001: out_v[16] = 10'b0111000001;
    default: out_v[16] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010000010000010: out_v[17] = 10'b0011100001;
    16'b0011010100000100: out_v[17] = 10'b0111000110;
    16'b0011010110010010: out_v[17] = 10'b1011001011;
    16'b0000000010010010: out_v[17] = 10'b0101100001;
    16'b0011010000000000: out_v[17] = 10'b1100110011;
    16'b0010000000000000: out_v[17] = 10'b1111000010;
    16'b0010010000000100: out_v[17] = 10'b1100011110;
    16'b0010000010010000: out_v[17] = 10'b0010001100;
    16'b0010010010000110: out_v[17] = 10'b1010101100;
    16'b0010000010010010: out_v[17] = 10'b0100111011;
    16'b0010000110000010: out_v[17] = 10'b1101010000;
    16'b0010000010000000: out_v[17] = 10'b1100100101;
    16'b0000000000000000: out_v[17] = 10'b1010000001;
    16'b0010010100100000: out_v[17] = 10'b0001001000;
    16'b0011010100000000: out_v[17] = 10'b0010101111;
    16'b0011010110110010: out_v[17] = 10'b1111100010;
    16'b0000000010000010: out_v[17] = 10'b1011000001;
    16'b0011010100100000: out_v[17] = 10'b1100001111;
    16'b0000000000000010: out_v[17] = 10'b0000011000;
    16'b0011010000000100: out_v[17] = 10'b0011011011;
    16'b0010010110110010: out_v[17] = 10'b0001101110;
    16'b0011010110100010: out_v[17] = 10'b1111000011;
    16'b0010000000000100: out_v[17] = 10'b0100100011;
    16'b0010000000000010: out_v[17] = 10'b0011000110;
    16'b0000000010010000: out_v[17] = 10'b0100100001;
    16'b0011000010010010: out_v[17] = 10'b0010001101;
    16'b0011010100100100: out_v[17] = 10'b1001010111;
    16'b0010010010010010: out_v[17] = 10'b0000000111;
    16'b0010000110010010: out_v[17] = 10'b0010100100;
    16'b0011010110110000: out_v[17] = 10'b1011110110;
    16'b0011010110100110: out_v[17] = 10'b1111110011;
    16'b0010010000000000: out_v[17] = 10'b1000010101;
    16'b0011010010010010: out_v[17] = 10'b0011000011;
    16'b0010000110000000: out_v[17] = 10'b0001001001;
    16'b0000000100100000: out_v[17] = 10'b0000110111;
    16'b0001010000000000: out_v[17] = 10'b0110011010;
    16'b0011010110100000: out_v[17] = 10'b1111010000;
    16'b0000000000010000: out_v[17] = 10'b0001110000;
    16'b0010000110010000: out_v[17] = 10'b1011011110;
    16'b0010000000010000: out_v[17] = 10'b0001001010;
    16'b0010010110010010: out_v[17] = 10'b1001111011;
    16'b0001010100100000: out_v[17] = 10'b0111101001;
    16'b0011010110110110: out_v[17] = 10'b1000010011;
    16'b0000000010000000: out_v[17] = 10'b0110110001;
    16'b0000000100000000: out_v[17] = 10'b0010100101;
    16'b0010010110110000: out_v[17] = 10'b1111001011;
    16'b0010000100100000: out_v[17] = 10'b0001011110;
    16'b0010010010010000: out_v[17] = 10'b1111000111;
    16'b0001000100100000: out_v[17] = 10'b0101100001;
    16'b0001000000000000: out_v[17] = 10'b1010100100;
    16'b0000000100110000: out_v[17] = 10'b1011101111;
    16'b0010000110110010: out_v[17] = 10'b0010100100;
    16'b0000010000000000: out_v[17] = 10'b0001011100;
    16'b0000000110110010: out_v[17] = 10'b1011001000;
    16'b0010000110110000: out_v[17] = 10'b0011111010;
    16'b0000010010010000: out_v[17] = 10'b0110110110;
    16'b0010010010000010: out_v[17] = 10'b0001000000;
    16'b0000000110110000: out_v[17] = 10'b0011011110;
    16'b0010000010110010: out_v[17] = 10'b1010001111;
    16'b0010000000010010: out_v[17] = 10'b1100011101;
    16'b0011000110110010: out_v[17] = 10'b0010100100;
    16'b0000010010010010: out_v[17] = 10'b1111100110;
    16'b0010000110100010: out_v[17] = 10'b0011011100;
    16'b0011000000000000: out_v[17] = 10'b1101111110;
    16'b0000000110100000: out_v[17] = 10'b0001111000;
    16'b0001000100000000: out_v[17] = 10'b1100100110;
    16'b0000010110100000: out_v[17] = 10'b1100010011;
    16'b0000010100100000: out_v[17] = 10'b1101001010;
    16'b0000000100101000: out_v[17] = 10'b1001100111;
    16'b0000000110000000: out_v[17] = 10'b1011100011;
    16'b0000000110010010: out_v[17] = 10'b0001100011;
    16'b0000000110000010: out_v[17] = 10'b1011101100;
    16'b0010000110100000: out_v[17] = 10'b1101001011;
    16'b0000010100000000: out_v[17] = 10'b1010001110;
    16'b0010000100000000: out_v[17] = 10'b1011010111;
    16'b0000000110100010: out_v[17] = 10'b1100100011;
    16'b0000000110010000: out_v[17] = 10'b0000010011;
    16'b0001000000000010: out_v[17] = 10'b0101110001;
    16'b0000010000000010: out_v[17] = 10'b1000110010;
    16'b0001000100101000: out_v[17] = 10'b1010010100;
    16'b0001000100000010: out_v[17] = 10'b0110111111;
    16'b0000000100000010: out_v[17] = 10'b1110100110;
    16'b0000000100100010: out_v[17] = 10'b0010101010;
    16'b0001000100100010: out_v[17] = 10'b0110001111;
    16'b0001000110101000: out_v[17] = 10'b0111001100;
    16'b0001000110100010: out_v[17] = 10'b1010101111;
    16'b0001000100101010: out_v[17] = 10'b1011000111;
    16'b0001010110110010: out_v[17] = 10'b1100100111;
    16'b0001010110100010: out_v[17] = 10'b0100100110;
    16'b0001010000000100: out_v[17] = 10'b0001100001;
    16'b0000010000010000: out_v[17] = 10'b0110111010;
    16'b0010010000010000: out_v[17] = 10'b1001111010;
    16'b0001010000010000: out_v[17] = 10'b1111011000;
    16'b0000000100010000: out_v[17] = 10'b0000110010;
    16'b0001000010000010: out_v[17] = 10'b0001011111;
    16'b0001000110100000: out_v[17] = 10'b0110001111;
    16'b0001000000101000: out_v[17] = 10'b1111001010;
    default: out_v[17] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1010000000010000: out_v[18] = 10'b0010001010;
    16'b0010000000011000: out_v[18] = 10'b1101010101;
    16'b1010110101101000: out_v[18] = 10'b0001111100;
    16'b1010110100001000: out_v[18] = 10'b1101111011;
    16'b1010000100010000: out_v[18] = 10'b0010110011;
    16'b0010000100010000: out_v[18] = 10'b0110100011;
    16'b1010110000101000: out_v[18] = 10'b1101110110;
    16'b1010010000101000: out_v[18] = 10'b1010001111;
    16'b0010000100111000: out_v[18] = 10'b0111111110;
    16'b1010010000011000: out_v[18] = 10'b0011000010;
    16'b1010010000000000: out_v[18] = 10'b0011100011;
    16'b1010010000001000: out_v[18] = 10'b0001011011;
    16'b1010000000001000: out_v[18] = 10'b1011101111;
    16'b1011110100101000: out_v[18] = 10'b1111111000;
    16'b1010110101001000: out_v[18] = 10'b1111111010;
    16'b1010010100001000: out_v[18] = 10'b0111110100;
    16'b0010000000010000: out_v[18] = 10'b0011010111;
    16'b1010000100011000: out_v[18] = 10'b1100010010;
    16'b1010010100000000: out_v[18] = 10'b1101110110;
    16'b0010000100011000: out_v[18] = 10'b1010001011;
    16'b1011110101101000: out_v[18] = 10'b1111100010;
    16'b1011110001101000: out_v[18] = 10'b0101000111;
    16'b1010110100111000: out_v[18] = 10'b1111010011;
    16'b1010110100101000: out_v[18] = 10'b1011110010;
    16'b1010110001101000: out_v[18] = 10'b1100001111;
    16'b1010010000010000: out_v[18] = 10'b0111110100;
    16'b1010010100011000: out_v[18] = 10'b1100111111;
    16'b1010000100001000: out_v[18] = 10'b1111000111;
    16'b1010000000000000: out_v[18] = 10'b0100001101;
    16'b1010000000011000: out_v[18] = 10'b0011001111;
    16'b1011110000101000: out_v[18] = 10'b1000101111;
    16'b1010110000001000: out_v[18] = 10'b0111111011;
    16'b1010000100111000: out_v[18] = 10'b0100100111;
    16'b1010010100010000: out_v[18] = 10'b1011110011;
    16'b1010010100101000: out_v[18] = 10'b1101110110;
    16'b1010000100010010: out_v[18] = 10'b1101001011;
    16'b1010010100111000: out_v[18] = 10'b1111010111;
    16'b0010000100000110: out_v[18] = 10'b0000100111;
    16'b0000000000000100: out_v[18] = 10'b0101001010;
    16'b0000000100000110: out_v[18] = 10'b1001110111;
    16'b0000000000000110: out_v[18] = 10'b1010101111;
    16'b0010000000000110: out_v[18] = 10'b1100100100;
    16'b1000000000000100: out_v[18] = 10'b1000000011;
    16'b1000000000000110: out_v[18] = 10'b0010001011;
    16'b0000000100000010: out_v[18] = 10'b1101000010;
    16'b0000000100000100: out_v[18] = 10'b0100011101;
    16'b0000000000000000: out_v[18] = 10'b0000011101;
    16'b1000000100000110: out_v[18] = 10'b0110000111;
    16'b0000000000000010: out_v[18] = 10'b0010111010;
    16'b0000001100000110: out_v[18] = 10'b1010000101;
    16'b0010001100010100: out_v[18] = 10'b1110110100;
    16'b1011000100000110: out_v[18] = 10'b1010111011;
    16'b0010001100000110: out_v[18] = 10'b0000111100;
    16'b1010000100000000: out_v[18] = 10'b1001110110;
    16'b0010000100000010: out_v[18] = 10'b1001001000;
    16'b0010001100000010: out_v[18] = 10'b1111011000;
    16'b1010000100001010: out_v[18] = 10'b1001011110;
    16'b1010000100000010: out_v[18] = 10'b0100001111;
    16'b1010000100000110: out_v[18] = 10'b0111010101;
    16'b1010001100000010: out_v[18] = 10'b1111001111;
    16'b1010010100000110: out_v[18] = 10'b0110000101;
    16'b1000000100000010: out_v[18] = 10'b0101110101;
    16'b1001010100000110: out_v[18] = 10'b1110001101;
    16'b1010001100000110: out_v[18] = 10'b0111100001;
    16'b0000001100000010: out_v[18] = 10'b0110101100;
    16'b0010000100000000: out_v[18] = 10'b0111000101;
    16'b1010000000000010: out_v[18] = 10'b1100101110;
    16'b1010010100000010: out_v[18] = 10'b0010110100;
    16'b0010001100010110: out_v[18] = 10'b0010110101;
    16'b1010000000000110: out_v[18] = 10'b0100010011;
    16'b0010000100001010: out_v[18] = 10'b1011001100;
    16'b0010000000000010: out_v[18] = 10'b1011101001;
    16'b0011001100000110: out_v[18] = 10'b1111111011;
    16'b1001000100000110: out_v[18] = 10'b1110111011;
    16'b0010001100010000: out_v[18] = 10'b1100100111;
    16'b0001000100000110: out_v[18] = 10'b0010011011;
    16'b0010001100010010: out_v[18] = 10'b0100101011;
    16'b0010001100000000: out_v[18] = 10'b1100001110;
    16'b1010010000010100: out_v[18] = 10'b1101001010;
    16'b0000000000010100: out_v[18] = 10'b0101011010;
    16'b0010000100000100: out_v[18] = 10'b1100001001;
    16'b1010000100000100: out_v[18] = 10'b1001001001;
    16'b1000000000010100: out_v[18] = 10'b0010110110;
    16'b1010000000010110: out_v[18] = 10'b1000111110;
    16'b0010000000000100: out_v[18] = 10'b1000011011;
    16'b0010000000010100: out_v[18] = 10'b1001101000;
    16'b1010000000010100: out_v[18] = 10'b0101110110;
    16'b0010000100010100: out_v[18] = 10'b1001101110;
    16'b1010000100010100: out_v[18] = 10'b0010111110;
    16'b1010000000000100: out_v[18] = 10'b1110010011;
    16'b0000000100010100: out_v[18] = 10'b0001001110;
    16'b1000010000000100: out_v[18] = 10'b0111001011;
    16'b1000000100000100: out_v[18] = 10'b0100111111;
    16'b0010001100000100: out_v[18] = 10'b1010011000;
    16'b0010000100011100: out_v[18] = 10'b0011101000;
    16'b1010000100011100: out_v[18] = 10'b0011101111;
    16'b1000000000000000: out_v[18] = 10'b1110100100;
    16'b1010010000000100: out_v[18] = 10'b1101101010;
    16'b1010000000001100: out_v[18] = 10'b1111001111;
    16'b1010010100010100: out_v[18] = 10'b1001101110;
    16'b0010000000000000: out_v[18] = 10'b0111001001;
    16'b0010010000000100: out_v[18] = 10'b0110011000;
    16'b1010000100001100: out_v[18] = 10'b1001011001;
    16'b1000000100010100: out_v[18] = 10'b1001001101;
    16'b1010010000000110: out_v[18] = 10'b0011011111;
    16'b1010010100000100: out_v[18] = 10'b1000101011;
    16'b0010010000010110: out_v[18] = 10'b0001101101;
    16'b0010000100010110: out_v[18] = 10'b1001011101;
    16'b0010010000010100: out_v[18] = 10'b0101100101;
    16'b0000000100010010: out_v[18] = 10'b1111000010;
    16'b1010000100010110: out_v[18] = 10'b0101110001;
    16'b1000000100010110: out_v[18] = 10'b0011101011;
    16'b1010010100010110: out_v[18] = 10'b1100010010;
    16'b1000000000010010: out_v[18] = 10'b1000111100;
    16'b1000000000010110: out_v[18] = 10'b1000111111;
    16'b1000010000010010: out_v[18] = 10'b1010001100;
    16'b1010000000010010: out_v[18] = 10'b1100110010;
    16'b1010010000010110: out_v[18] = 10'b1010110010;
    16'b0010110001000010: out_v[18] = 10'b0111111011;
    16'b1000000000000010: out_v[18] = 10'b1000011100;
    16'b0010010000000010: out_v[18] = 10'b0111110110;
    16'b0010010000010000: out_v[18] = 10'b0111101110;
    16'b0010000000010010: out_v[18] = 10'b1001001010;
    16'b1000010000010100: out_v[18] = 10'b1100000101;
    16'b0000000100010110: out_v[18] = 10'b0001010001;
    16'b0000010000010100: out_v[18] = 10'b0000111000;
    16'b0010010000010010: out_v[18] = 10'b1011110011;
    16'b1010010000010010: out_v[18] = 10'b1000111110;
    16'b0000010000000010: out_v[18] = 10'b0000011110;
    16'b0010000000010110: out_v[18] = 10'b1001001101;
    16'b0000110001001010: out_v[18] = 10'b1101111101;
    16'b0000000000010110: out_v[18] = 10'b1100111100;
    16'b0000000000010010: out_v[18] = 10'b0101111110;
    16'b1000000000010000: out_v[18] = 10'b0010000111;
    16'b0010010000000110: out_v[18] = 10'b0110010011;
    16'b0010110001010100: out_v[18] = 10'b0000111100;
    16'b1010010000000010: out_v[18] = 10'b1101101110;
    16'b1000010000000010: out_v[18] = 10'b1100101010;
    16'b1000110000001010: out_v[18] = 10'b1110010001;
    16'b0000000100011000: out_v[18] = 10'b0000001011;
    16'b0010000100010010: out_v[18] = 10'b1001000100;
    16'b0000000100011100: out_v[18] = 10'b0011110011;
    16'b0000000100010000: out_v[18] = 10'b1111000010;
    16'b0000000100001100: out_v[18] = 10'b0101110101;
    16'b0000000100011010: out_v[18] = 10'b1100101010;
    16'b1000000100010000: out_v[18] = 10'b1100100011;
    16'b1000000100010010: out_v[18] = 10'b0000001011;
    16'b1000001100010110: out_v[18] = 10'b1010000101;
    16'b1000001100010100: out_v[18] = 10'b1111000110;
    16'b1000011100010110: out_v[18] = 10'b0001001110;
    16'b1000001100010010: out_v[18] = 10'b0111100010;
    16'b1000001100010000: out_v[18] = 10'b1111001000;
    16'b1000001100000110: out_v[18] = 10'b1001010011;
    16'b1000011100010010: out_v[18] = 10'b1011001000;
    16'b0000001100010010: out_v[18] = 10'b1111101010;
    16'b1000010100010110: out_v[18] = 10'b0111001011;
    16'b0000001100010110: out_v[18] = 10'b1101101001;
    16'b1000001100000010: out_v[18] = 10'b1100011011;
    16'b1000011100000110: out_v[18] = 10'b0011101011;
    16'b1000011100000000: out_v[18] = 10'b0110001111;
    16'b1000010100000110: out_v[18] = 10'b0010100011;
    16'b1000011100000100: out_v[18] = 10'b1000110011;
    16'b1010010101001000: out_v[18] = 10'b0111010110;
    16'b1000010001000000: out_v[18] = 10'b1111110111;
    16'b1000010000000000: out_v[18] = 10'b1001100010;
    16'b1000010100000000: out_v[18] = 10'b0111110000;
    16'b0000010000000000: out_v[18] = 10'b0011110100;
    16'b1010010001000100: out_v[18] = 10'b0011111111;
    16'b1010000100001110: out_v[18] = 10'b0111110011;
    16'b1010010001000000: out_v[18] = 10'b1011010011;
    16'b1000010000010000: out_v[18] = 10'b0010101110;
    16'b1010010101000000: out_v[18] = 10'b0101111110;
    16'b1000000100000000: out_v[18] = 10'b0111100000;
    16'b0000010001000000: out_v[18] = 10'b0011010001;
    16'b1000010100001000: out_v[18] = 10'b1001011100;
    16'b1000010001001000: out_v[18] = 10'b0001011110;
    16'b1010010101000100: out_v[18] = 10'b0010111001;
    16'b1000010000001000: out_v[18] = 10'b0011111111;
    16'b1000010101001000: out_v[18] = 10'b1101011011;
    16'b1010010100001110: out_v[18] = 10'b1101000001;
    16'b1000010000000110: out_v[18] = 10'b0010101010;
    16'b1010110001000000: out_v[18] = 10'b0110101111;
    16'b1000010001000100: out_v[18] = 10'b0111110001;
    16'b1010010100001010: out_v[18] = 10'b1100000111;
    16'b1010000000011110: out_v[18] = 10'b0001011011;
    16'b0010000100001110: out_v[18] = 10'b1110100000;
    16'b1010010100011110: out_v[18] = 10'b0110100011;
    16'b0010000000001110: out_v[18] = 10'b1111010101;
    16'b1010010101010110: out_v[18] = 10'b0101100100;
    16'b1010000000001110: out_v[18] = 10'b0101000011;
    16'b1010010000001110: out_v[18] = 10'b0001000111;
    16'b1000000000001110: out_v[18] = 10'b1110000011;
    16'b0010010100000110: out_v[18] = 10'b1110010001;
    16'b1010010000011110: out_v[18] = 10'b0111110100;
    16'b1010000100011110: out_v[18] = 10'b1010100011;
    16'b0000010100000110: out_v[18] = 10'b1110000101;
    16'b1010110001001010: out_v[18] = 10'b1101001011;
    16'b1010110001000010: out_v[18] = 10'b1101001011;
    16'b1010010100011100: out_v[18] = 10'b1001101010;
    16'b1010110001000110: out_v[18] = 10'b1101110111;
    16'b1000110001000010: out_v[18] = 10'b1000000010;
    16'b1000010000010110: out_v[18] = 10'b1100100111;
    default: out_v[18] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0101100101000000: out_v[19] = 10'b0110011001;
    16'b0101101100000001: out_v[19] = 10'b0000110101;
    16'b0001101101100011: out_v[19] = 10'b0111110001;
    16'b0101101100000000: out_v[19] = 10'b1100010010;
    16'b0001101001000011: out_v[19] = 10'b1000001011;
    16'b0001101000000001: out_v[19] = 10'b1100001101;
    16'b0101101101000001: out_v[19] = 10'b0111010100;
    16'b0101101101000000: out_v[19] = 10'b0000001011;
    16'b0101101101000011: out_v[19] = 10'b1100000111;
    16'b0001001101000001: out_v[19] = 10'b0000001011;
    16'b0101100001000000: out_v[19] = 10'b1010100111;
    16'b0001101001000010: out_v[19] = 10'b1110101011;
    16'b0101101001000001: out_v[19] = 10'b0010101110;
    16'b0101001101000001: out_v[19] = 10'b1001001110;
    16'b0101101101100011: out_v[19] = 10'b1010100111;
    16'b0100001101000001: out_v[19] = 10'b0110001111;
    16'b0001101000000011: out_v[19] = 10'b1001111010;
    16'b0001101101000011: out_v[19] = 10'b1110111010;
    16'b0001101101000001: out_v[19] = 10'b1100110100;
    16'b0001101101000000: out_v[19] = 10'b1001011100;
    16'b0101101001000011: out_v[19] = 10'b1100000001;
    16'b0001101101001011: out_v[19] = 10'b1011010011;
    16'b0001101001000001: out_v[19] = 10'b0111110111;
    16'b0101101000000001: out_v[19] = 10'b1010001111;
    16'b0101101111000001: out_v[19] = 10'b1010011111;
    16'b0001101100000011: out_v[19] = 10'b1100011101;
    16'b0001101001001011: out_v[19] = 10'b1110010111;
    16'b0000001101000001: out_v[19] = 10'b0111000011;
    16'b0101101001100011: out_v[19] = 10'b1000000011;
    16'b0101100100000000: out_v[19] = 10'b0110011000;
    16'b0001101001100011: out_v[19] = 10'b0111111111;
    16'b0101101001000000: out_v[19] = 10'b0110111010;
    16'b0101101101100001: out_v[19] = 10'b1011001111;
    16'b0001100101100011: out_v[19] = 10'b1011110010;
    16'b0101101000000000: out_v[19] = 10'b0100010101;
    16'b0000001100000001: out_v[19] = 10'b1100000001;
    16'b0101100101000001: out_v[19] = 10'b0001011011;
    16'b0101001101000011: out_v[19] = 10'b0110110110;
    16'b0001100001100011: out_v[19] = 10'b0111110001;
    16'b0001001101000011: out_v[19] = 10'b1110111110;
    16'b0101101110000001: out_v[19] = 10'b0010011011;
    16'b0001101001000000: out_v[19] = 10'b1110100111;
    16'b0001100100000000: out_v[19] = 10'b0001011011;
    16'b0001000001000000: out_v[19] = 10'b1010000011;
    16'b0000000001000000: out_v[19] = 10'b0000011011;
    16'b0001000000000000: out_v[19] = 10'b0010011001;
    16'b0000000000000000: out_v[19] = 10'b0110111111;
    16'b0000100000000000: out_v[19] = 10'b1110100001;
    16'b0001100000000000: out_v[19] = 10'b0111010001;
    16'b0000100010000000: out_v[19] = 10'b1011100110;
    16'b0001000100000000: out_v[19] = 10'b1111001001;
    16'b0001100001000000: out_v[19] = 10'b1001101000;
    16'b0001100010000000: out_v[19] = 10'b0010101110;
    16'b0001100101000000: out_v[19] = 10'b1000010010;
    16'b0000100100000000: out_v[19] = 10'b0110010011;
    16'b0001000101000000: out_v[19] = 10'b0101110101;
    16'b0001100001001000: out_v[19] = 10'b0101000110;
    16'b0000101100000000: out_v[19] = 10'b1110001101;
    16'b0001101100000000: out_v[19] = 10'b0000010111;
    16'b0101100000000000: out_v[19] = 10'b0110110100;
    16'b0001100000001000: out_v[19] = 10'b0001011100;
    16'b0100101100000000: out_v[19] = 10'b1100001110;
    16'b0100001100100001: out_v[19] = 10'b1010111110;
    16'b0000000100000000: out_v[19] = 10'b1111001000;
    16'b0001101000000000: out_v[19] = 10'b1100000110;
    16'b0001101101001000: out_v[19] = 10'b0010110110;
    16'b0100001100000000: out_v[19] = 10'b1010110110;
    16'b0000101101000000: out_v[19] = 10'b1001010111;
    16'b0000001101000000: out_v[19] = 10'b1111001110;
    16'b0001001101000000: out_v[19] = 10'b0011101010;
    16'b0001100101001000: out_v[19] = 10'b1100001100;
    16'b0100001001000000: out_v[19] = 10'b0111011001;
    16'b0000100101000000: out_v[19] = 10'b1110100000;
    16'b0000001001000000: out_v[19] = 10'b0100010101;
    16'b0100001100000001: out_v[19] = 10'b0101000110;
    16'b0001100100001000: out_v[19] = 10'b0000011010;
    16'b0100000001000000: out_v[19] = 10'b0001011110;
    16'b0000001100000000: out_v[19] = 10'b1111100101;
    16'b0100100101000000: out_v[19] = 10'b1101001011;
    16'b0001100001000001: out_v[19] = 10'b1000101010;
    16'b0101000101000000: out_v[19] = 10'b0010100110;
    16'b0101000001000000: out_v[19] = 10'b1001011101;
    16'b0101100001001000: out_v[19] = 10'b1010100000;
    16'b0001000101000001: out_v[19] = 10'b0001111110;
    16'b0101100000001000: out_v[19] = 10'b0111011110;
    16'b0101000001001000: out_v[19] = 10'b1101100101;
    16'b0101100101001000: out_v[19] = 10'b0001001010;
    16'b0100000100000000: out_v[19] = 10'b0001100001;
    16'b0101100001000001: out_v[19] = 10'b1111001010;
    16'b0100100100000000: out_v[19] = 10'b1100001101;
    16'b0100000001001000: out_v[19] = 10'b1001001101;
    16'b0101000101000001: out_v[19] = 10'b1100001011;
    16'b0101000000000000: out_v[19] = 10'b0100011000;
    16'b0001100101000001: out_v[19] = 10'b0001111000;
    16'b0000000001000001: out_v[19] = 10'b0011110111;
    16'b0100100000000000: out_v[19] = 10'b0110001010;
    16'b0100000001000001: out_v[19] = 10'b0001011111;
    16'b0100000000000001: out_v[19] = 10'b1000101001;
    16'b0100100001000000: out_v[19] = 10'b0010010111;
    16'b0100100000000010: out_v[19] = 10'b0100001001;
    16'b0100001001000001: out_v[19] = 10'b0111111000;
    16'b0100000000000011: out_v[19] = 10'b0111001110;
    16'b0000001010000000: out_v[19] = 10'b1011011101;
    16'b0000101000000000: out_v[19] = 10'b1101100110;
    16'b0100000000001000: out_v[19] = 10'b0010011100;
    16'b0100000000000000: out_v[19] = 10'b0011100111;
    16'b0100001000000001: out_v[19] = 10'b1001011010;
    16'b0101101100001010: out_v[19] = 10'b0101011000;
    16'b0100001000000010: out_v[19] = 10'b1001011011;
    16'b0100101000000000: out_v[19] = 10'b1111001101;
    16'b0000001000000000: out_v[19] = 10'b0001101110;
    16'b0000100001000000: out_v[19] = 10'b0001111101;
    16'b0100001010000000: out_v[19] = 10'b1111100010;
    16'b0100000000000010: out_v[19] = 10'b0110100101;
    16'b0100001000000000: out_v[19] = 10'b0110000111;
    16'b0100001000001011: out_v[19] = 10'b0010111001;
    16'b0100101001000000: out_v[19] = 10'b0100011011;
    16'b0100001000000011: out_v[19] = 10'b0010011111;
    16'b0101100000001010: out_v[19] = 10'b0100010110;
    16'b0000001000000001: out_v[19] = 10'b1010101011;
    16'b0101100100001010: out_v[19] = 10'b0111011011;
    16'b0100100000001000: out_v[19] = 10'b0111110010;
    16'b0100000001000011: out_v[19] = 10'b0101010011;
    16'b0000000000000001: out_v[19] = 10'b0010100110;
    16'b0100001000100011: out_v[19] = 10'b0110111011;
    16'b0101100101000010: out_v[19] = 10'b0011101010;
    16'b0101000111000000: out_v[19] = 10'b1111100001;
    16'b0101100111000000: out_v[19] = 10'b0111000001;
    16'b0100000101000000: out_v[19] = 10'b1111100110;
    16'b0101100001000010: out_v[19] = 10'b1100100110;
    16'b0101000101001000: out_v[19] = 10'b0010101101;
    16'b0001100111000000: out_v[19] = 10'b1100111011;
    16'b0101100001001010: out_v[19] = 10'b0111100110;
    16'b0000101000000001: out_v[19] = 10'b1101011010;
    16'b0000000101000000: out_v[19] = 10'b1100100101;
    16'b0000100000000001: out_v[19] = 10'b1011110100;
    16'b0101100101001010: out_v[19] = 10'b0110110010;
    16'b0001100000000001: out_v[19] = 10'b1101001100;
    16'b0101001101000000: out_v[19] = 10'b1011100110;
    16'b0101000100000000: out_v[19] = 10'b1001011001;
    16'b0110000000000000: out_v[19] = 10'b1011000011;
    16'b0000001000000011: out_v[19] = 10'b0011010000;
    16'b0010000000000000: out_v[19] = 10'b0011000011;
    16'b0100001101000000: out_v[19] = 10'b1111000111;
    16'b0100001001000010: out_v[19] = 10'b1011100001;
    16'b0101101010000000: out_v[19] = 10'b0011000010;
    16'b0110001000000010: out_v[19] = 10'b1011111011;
    16'b0000001000000010: out_v[19] = 10'b0011001011;
    16'b0101001100000000: out_v[19] = 10'b1101100011;
    16'b0101101110000000: out_v[19] = 10'b1111010010;
    16'b0001100110000000: out_v[19] = 10'b1000110001;
    16'b0101100000000011: out_v[19] = 10'b0110010101;
    16'b0000100000000010: out_v[19] = 10'b0000110111;
    16'b0001100000000010: out_v[19] = 10'b0111110001;
    16'b0000100000000011: out_v[19] = 10'b1101101111;
    16'b0000100001000001: out_v[19] = 10'b1101100010;
    16'b0101100000000001: out_v[19] = 10'b1101011010;
    16'b0100100000000001: out_v[19] = 10'b1001011100;
    16'b0100100000000011: out_v[19] = 10'b0011110000;
    16'b0101100001000011: out_v[19] = 10'b1001100100;
    16'b0001100001000010: out_v[19] = 10'b0001101100;
    16'b0101100000000010: out_v[19] = 10'b1101011110;
    16'b0000000100000001: out_v[19] = 10'b1110001111;
    16'b0001000100000001: out_v[19] = 10'b1110101100;
    16'b0001100001000011: out_v[19] = 10'b1100100010;
    16'b0001000001000001: out_v[19] = 10'b1101100011;
    16'b0000000101000001: out_v[19] = 10'b1110001001;
    16'b0001100100000001: out_v[19] = 10'b0111110001;
    16'b0101101001001010: out_v[19] = 10'b1011101010;
    16'b0101100001011010: out_v[19] = 10'b1010001111;
    16'b0101101001000010: out_v[19] = 10'b1111110111;
    16'b0001100001001010: out_v[19] = 10'b0110101001;
    16'b0101101001011010: out_v[19] = 10'b1101101110;
    default: out_v[19] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100001100001000: out_v[20] = 10'b0001110001;
    16'b0101011110000000: out_v[20] = 10'b1101011010;
    16'b0000011110001000: out_v[20] = 10'b0010111110;
    16'b0100011100001000: out_v[20] = 10'b1011100011;
    16'b0100001100000000: out_v[20] = 10'b0011001000;
    16'b0000011110000000: out_v[20] = 10'b0001010111;
    16'b0100011110000000: out_v[20] = 10'b0100100000;
    16'b0000001110000000: out_v[20] = 10'b1000001011;
    16'b0100011110001000: out_v[20] = 10'b0111111011;
    16'b0100011110000100: out_v[20] = 10'b0111111010;
    16'b0101011110001000: out_v[20] = 10'b1011011000;
    16'b0100011100000000: out_v[20] = 10'b0110100011;
    16'b0100010110001000: out_v[20] = 10'b0010011011;
    16'b0000011110101000: out_v[20] = 10'b1011101100;
    16'b0000001110000100: out_v[20] = 10'b0101100111;
    16'b0000011010101000: out_v[20] = 10'b1111110011;
    16'b0000011010000000: out_v[20] = 10'b0110010101;
    16'b0000011010001000: out_v[20] = 10'b0100010111;
    16'b0000010010001000: out_v[20] = 10'b0000000110;
    16'b0000010000001000: out_v[20] = 10'b1111010000;
    16'b0100011110001100: out_v[20] = 10'b1110101101;
    16'b0000000010001000: out_v[20] = 10'b1111000011;
    16'b0100010110000000: out_v[20] = 10'b1001110011;
    16'b0000011110100000: out_v[20] = 10'b1001011010;
    16'b0101011110000100: out_v[20] = 10'b0111111111;
    16'b0001011110001000: out_v[20] = 10'b0010110101;
    16'b0100010010000000: out_v[20] = 10'b0000110011;
    16'b0100001101001000: out_v[20] = 10'b0000110001;
    16'b0100000100001000: out_v[20] = 10'b0001111001;
    16'b0000011110001100: out_v[20] = 10'b1110111110;
    16'b0000011100001000: out_v[20] = 10'b0111011110;
    16'b0000011110000100: out_v[20] = 10'b0000011111;
    16'b0100010100001000: out_v[20] = 10'b1000101110;
    16'b0101011110001100: out_v[20] = 10'b0110110001;
    16'b0000001010001000: out_v[20] = 10'b1111010111;
    16'b0000010110001000: out_v[20] = 10'b1000110001;
    16'b0000000001000010: out_v[20] = 10'b1000111011;
    16'b0000001001000010: out_v[20] = 10'b0010100100;
    16'b0000001000001010: out_v[20] = 10'b1101110101;
    16'b0000000000000010: out_v[20] = 10'b1100110011;
    16'b0000001001001010: out_v[20] = 10'b1101100010;
    16'b0000001000001000: out_v[20] = 10'b1111000111;
    16'b0001000001000010: out_v[20] = 10'b0000100110;
    16'b0000000001001010: out_v[20] = 10'b1010101001;
    16'b0000001000000010: out_v[20] = 10'b0101101100;
    16'b0000001101000010: out_v[20] = 10'b1110000000;
    16'b0000000000000000: out_v[20] = 10'b0001110101;
    16'b0000001101001010: out_v[20] = 10'b1010010011;
    16'b0000001000000000: out_v[20] = 10'b1010000110;
    16'b0000000000001010: out_v[20] = 10'b1011111011;
    16'b0000001100001000: out_v[20] = 10'b0100011111;
    16'b0000000000001000: out_v[20] = 10'b1000001100;
    16'b0000001100000000: out_v[20] = 10'b1001001110;
    16'b0000001100001010: out_v[20] = 10'b0110011010;
    16'b0000000001001000: out_v[20] = 10'b1010100100;
    16'b0100000000001000: out_v[20] = 10'b0100001100;
    16'b0000001101000000: out_v[20] = 10'b0011011011;
    16'b0000001001001000: out_v[20] = 10'b1100110101;
    16'b0000011000001000: out_v[20] = 10'b0001001010;
    16'b0000001101001000: out_v[20] = 10'b1000001100;
    16'b0000001001000000: out_v[20] = 10'b0110100000;
    16'b0000000001000000: out_v[20] = 10'b0000010101;
    16'b0100000001001000: out_v[20] = 10'b1110100011;
    16'b0100000001001010: out_v[20] = 10'b1010001100;
    16'b0100001001001010: out_v[20] = 10'b0010001000;
    16'b0000000101001010: out_v[20] = 10'b0100000001;
    16'b0101000001001010: out_v[20] = 10'b1001000111;
    16'b0001001101001010: out_v[20] = 10'b1100001111;
    16'b0001001001000010: out_v[20] = 10'b0101011001;
    16'b0100010001001010: out_v[20] = 10'b1111101001;
    16'b0100001001000010: out_v[20] = 10'b1100100010;
    16'b0100001101001010: out_v[20] = 10'b1001000110;
    16'b0001000001001010: out_v[20] = 10'b0110101001;
    16'b0100000101001010: out_v[20] = 10'b1100010100;
    16'b0001001001001010: out_v[20] = 10'b1010110000;
    16'b0100001000000000: out_v[20] = 10'b1000101111;
    16'b0001000000001000: out_v[20] = 10'b1101011111;
    16'b0101001001000010: out_v[20] = 10'b0100001111;
    16'b0100011101001010: out_v[20] = 10'b0011101010;
    16'b0000010001001010: out_v[20] = 10'b1011001001;
    16'b0101001001001010: out_v[20] = 10'b0011011001;
    16'b0100011001001010: out_v[20] = 10'b0100010100;
    16'b0001001101000010: out_v[20] = 10'b1001111101;
    16'b0101001101001010: out_v[20] = 10'b0100010010;
    16'b0100001101000010: out_v[20] = 10'b1000001010;
    16'b0100000101001000: out_v[20] = 10'b0000001100;
    16'b0100000101000010: out_v[20] = 10'b0001010101;
    16'b0100000001000000: out_v[20] = 10'b1101110000;
    16'b0000000101000010: out_v[20] = 10'b1100000110;
    16'b0100000000000000: out_v[20] = 10'b1111110011;
    16'b0101001101000010: out_v[20] = 10'b1000000100;
    16'b0100000001000010: out_v[20] = 10'b0101010100;
    16'b0100001101000000: out_v[20] = 10'b0011001010;
    16'b0100000101000000: out_v[20] = 10'b0111010001;
    16'b0100010101000000: out_v[20] = 10'b0100111111;
    16'b0000000100000000: out_v[20] = 10'b0110100010;
    16'b0000010001000000: out_v[20] = 10'b1101110110;
    16'b0100011111000010: out_v[20] = 10'b0011111110;
    16'b0100010101000010: out_v[20] = 10'b1001001011;
    16'b0100011101000000: out_v[20] = 10'b1001011111;
    16'b0101001101000000: out_v[20] = 10'b0110110000;
    16'b0100010111000000: out_v[20] = 10'b1011110000;
    16'b0100011111000000: out_v[20] = 10'b1111110001;
    16'b0000010000000000: out_v[20] = 10'b0110000011;
    16'b0000000101000000: out_v[20] = 10'b0110000000;
    16'b0000010011000000: out_v[20] = 10'b1101111010;
    16'b0100010011000010: out_v[20] = 10'b0001010110;
    16'b0100001001000000: out_v[20] = 10'b1101110101;
    16'b0100011101000010: out_v[20] = 10'b1001100110;
    16'b0000010010000000: out_v[20] = 10'b0000011110;
    16'b0100010111000010: out_v[20] = 10'b0000111111;
    16'b0100010001000010: out_v[20] = 10'b0001010010;
    16'b0100000100000000: out_v[20] = 10'b0111001011;
    16'b0001001100000000: out_v[20] = 10'b0001011111;
    16'b0101001100000000: out_v[20] = 10'b0110100011;
    16'b0101001100001000: out_v[20] = 10'b1000100011;
    16'b0100011101001000: out_v[20] = 10'b0011010011;
    16'b0000010011010010: out_v[20] = 10'b1111111101;
    16'b0100011111001010: out_v[20] = 10'b0111011011;
    16'b0100011111001000: out_v[20] = 10'b1000110001;
    16'b0000010011001000: out_v[20] = 10'b1001001011;
    16'b0000010011001010: out_v[20] = 10'b1011111110;
    16'b0000010011000010: out_v[20] = 10'b0001001101;
    16'b0000011111001010: out_v[20] = 10'b0001010011;
    16'b0000011100000000: out_v[20] = 10'b1011001010;
    16'b0001001101000000: out_v[20] = 10'b0101011110;
    16'b0001001001000000: out_v[20] = 10'b0110111001;
    16'b0011001101000000: out_v[20] = 10'b0101010111;
    16'b0000011101000010: out_v[20] = 10'b1011101010;
    16'b0000001101100000: out_v[20] = 10'b0010111111;
    16'b0000001100100000: out_v[20] = 10'b0001110110;
    16'b0001001101001000: out_v[20] = 10'b0001110011;
    16'b0000000101001000: out_v[20] = 10'b1100110000;
    16'b0100001001001000: out_v[20] = 10'b0110010111;
    16'b0000000100001000: out_v[20] = 10'b1100110101;
    default: out_v[20] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000000000000: out_v[21] = 10'b1010100011;
    16'b0000000001000110: out_v[21] = 10'b1000000101;
    16'b0000000001000101: out_v[21] = 10'b1110000101;
    16'b0000000000000100: out_v[21] = 10'b1001011100;
    16'b0000000001000100: out_v[21] = 10'b1010010001;
    16'b0000000100000100: out_v[21] = 10'b0110010110;
    16'b0000000001000000: out_v[21] = 10'b1010110011;
    16'b0000000000000110: out_v[21] = 10'b0000101010;
    16'b1000000001000000: out_v[21] = 10'b0100110011;
    16'b1000000001000100: out_v[21] = 10'b1011100111;
    16'b0000000001000111: out_v[21] = 10'b0010000101;
    16'b0000000001000001: out_v[21] = 10'b1110000111;
    16'b0000000101000110: out_v[21] = 10'b0000011110;
    16'b0000000001000011: out_v[21] = 10'b0111000011;
    16'b0000000001000010: out_v[21] = 10'b0111110011;
    16'b0000000101000101: out_v[21] = 10'b0110001100;
    16'b0000000101000100: out_v[21] = 10'b0101010100;
    16'b0000000100000000: out_v[21] = 10'b1011000100;
    16'b0000000000000010: out_v[21] = 10'b0011101100;
    16'b0000000100000010: out_v[21] = 10'b1011010011;
    16'b1000000100000000: out_v[21] = 10'b0000111001;
    16'b1001000100000100: out_v[21] = 10'b0100000101;
    16'b0001000000000100: out_v[21] = 10'b0011011001;
    16'b1001000000000100: out_v[21] = 10'b0000011101;
    16'b1000000000000100: out_v[21] = 10'b0001011110;
    16'b0001000100000100: out_v[21] = 10'b1011100100;
    16'b1000000100000100: out_v[21] = 10'b1110000100;
    16'b0000000101000000: out_v[21] = 10'b1101110101;
    16'b1000000000000000: out_v[21] = 10'b0100110000;
    16'b1001000100000000: out_v[21] = 10'b0010111001;
    16'b0000000100000110: out_v[21] = 10'b0100101100;
    16'b0001000100000000: out_v[21] = 10'b0010011100;
    16'b1000000100000110: out_v[21] = 10'b1110100011;
    16'b0000001100000100: out_v[21] = 10'b1100000011;
    16'b0001001100000100: out_v[21] = 10'b0011100111;
    16'b1000000101000100: out_v[21] = 10'b0111000111;
    16'b1000000000000010: out_v[21] = 10'b1010101100;
    16'b1000000000000110: out_v[21] = 10'b1000111000;
    16'b0000000100100000: out_v[21] = 10'b0010011100;
    16'b0000000000100000: out_v[21] = 10'b0101101111;
    16'b1000010000000000: out_v[21] = 10'b1100011000;
    16'b0000000100100100: out_v[21] = 10'b1100000010;
    16'b1000000100000010: out_v[21] = 10'b0011011001;
    16'b0010000100000000: out_v[21] = 10'b1111101101;
    16'b0010000000000000: out_v[21] = 10'b1011111100;
    16'b0100000100000001: out_v[21] = 10'b1011111101;
    16'b0100000100000101: out_v[21] = 10'b0010101110;
    16'b0010000000000100: out_v[21] = 10'b0110110010;
    16'b0100000100000000: out_v[21] = 10'b1001101111;
    16'b0010000100000100: out_v[21] = 10'b1001101000;
    16'b0100000000000100: out_v[21] = 10'b0011101100;
    16'b0010000100000110: out_v[21] = 10'b1111000011;
    16'b0100000000000000: out_v[21] = 10'b1001111110;
    16'b0100000100000100: out_v[21] = 10'b0111101111;
    16'b0000000100000001: out_v[21] = 10'b1111100010;
    16'b0000000100000101: out_v[21] = 10'b1011100010;
    16'b1001000101000100: out_v[21] = 10'b0011000110;
    16'b0000001000000100: out_v[21] = 10'b0011001010;
    16'b1001000001000100: out_v[21] = 10'b0110001001;
    16'b0001000101000100: out_v[21] = 10'b1111100001;
    16'b0000001101000100: out_v[21] = 10'b1011101000;
    16'b0001001101000100: out_v[21] = 10'b1101011101;
    16'b0001001001000100: out_v[21] = 10'b0111110111;
    16'b0001000001000100: out_v[21] = 10'b0111000010;
    16'b0000001001000100: out_v[21] = 10'b1101110100;
    16'b0000000000100100: out_v[21] = 10'b1111000110;
    16'b0000010100100100: out_v[21] = 10'b0011011001;
    16'b0000010100000100: out_v[21] = 10'b0011001111;
    16'b0000010000000100: out_v[21] = 10'b1010001001;
    16'b0000010000100100: out_v[21] = 10'b1010101110;
    16'b0000010000000000: out_v[21] = 10'b0111011010;
    16'b0000000001100100: out_v[21] = 10'b1111001110;
    16'b0100000101000101: out_v[21] = 10'b0100011100;
    16'b0000000101000011: out_v[21] = 10'b0110000110;
    16'b0000000101000001: out_v[21] = 10'b0100011111;
    16'b0000000101000010: out_v[21] = 10'b0110111001;
    16'b0000000101000111: out_v[21] = 10'b1110011011;
    16'b0000000101100100: out_v[21] = 10'b1010000011;
    default: out_v[21] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000010010000100: out_v[22] = 10'b0111010111;
    16'b0000010000001100: out_v[22] = 10'b0011010111;
    16'b0000010010001100: out_v[22] = 10'b0000101000;
    16'b0000010000001000: out_v[22] = 10'b1001001111;
    16'b0000010000000000: out_v[22] = 10'b0010001001;
    16'b0000010000010000: out_v[22] = 10'b0011000011;
    16'b0000000000000000: out_v[22] = 10'b0010100101;
    16'b0100010100000000: out_v[22] = 10'b1001111010;
    16'b0000010000011100: out_v[22] = 10'b1000000111;
    16'b0000000010001100: out_v[22] = 10'b1101110011;
    16'b0000010000011000: out_v[22] = 10'b0101100111;
    16'b0000000010000100: out_v[22] = 10'b0001110101;
    16'b0000110000010000: out_v[22] = 10'b1001010100;
    16'b0000010000000100: out_v[22] = 10'b1111011110;
    16'b0010000000000000: out_v[22] = 10'b1000110101;
    16'b0000000000010000: out_v[22] = 10'b0111001101;
    16'b0000010000000010: out_v[22] = 10'b1110100001;
    16'b0000010010010100: out_v[22] = 10'b0011100011;
    16'b0100100100011000: out_v[22] = 10'b1001100010;
    16'b0100100100010000: out_v[22] = 10'b0000110111;
    16'b0100100110000000: out_v[22] = 10'b1111000100;
    16'b0100100110000100: out_v[22] = 10'b0110000111;
    16'b0100100100000000: out_v[22] = 10'b1110101010;
    16'b0100100100001000: out_v[22] = 10'b0011011111;
    16'b0100000100010000: out_v[22] = 10'b0100010100;
    16'b0100110100010000: out_v[22] = 10'b0111100000;
    16'b0100100100010100: out_v[22] = 10'b1001010111;
    16'b0100100110010000: out_v[22] = 10'b1010000011;
    16'b0100000100000000: out_v[22] = 10'b0001010110;
    16'b0100100110010100: out_v[22] = 10'b0010010110;
    16'b0100100100000100: out_v[22] = 10'b1010010011;
    16'b0100110110010000: out_v[22] = 10'b0110010010;
    16'b0100010100010000: out_v[22] = 10'b0010111000;
    16'b0100000110000000: out_v[22] = 10'b1001011111;
    16'b0100000110010000: out_v[22] = 10'b1101010001;
    16'b0100110100000000: out_v[22] = 10'b0001000111;
    16'b0100100000000000: out_v[22] = 10'b1110001110;
    16'b0110110100010000: out_v[22] = 10'b0101010111;
    16'b0100100000011000: out_v[22] = 10'b1010110011;
    16'b0000100000010000: out_v[22] = 10'b0010011101;
    16'b0100110100001000: out_v[22] = 10'b1001111101;
    16'b0100110000010010: out_v[22] = 10'b0011100111;
    16'b0110110100000000: out_v[22] = 10'b0111001101;
    16'b0100110000010000: out_v[22] = 10'b0011001101;
    16'b0100010000010000: out_v[22] = 10'b0100011110;
    16'b0100100000010000: out_v[22] = 10'b0110010100;
    16'b0000110000011000: out_v[22] = 10'b1010011101;
    16'b0000110000010010: out_v[22] = 10'b1010101100;
    16'b0100110100010010: out_v[22] = 10'b1001000110;
    16'b0100000000010000: out_v[22] = 10'b0000101010;
    16'b0010110000010000: out_v[22] = 10'b0001001110;
    16'b0110100000010000: out_v[22] = 10'b1001011011;
    16'b0110100100010000: out_v[22] = 10'b0110000101;
    16'b0000110000000000: out_v[22] = 10'b0011101001;
    16'b0110110000010000: out_v[22] = 10'b0001000101;
    16'b0000100000010010: out_v[22] = 10'b0101000100;
    16'b0100110000011000: out_v[22] = 10'b1011101111;
    16'b0100110000000000: out_v[22] = 10'b0001001000;
    16'b0110010100000000: out_v[22] = 10'b0111000110;
    16'b0000100000011000: out_v[22] = 10'b0110010000;
    16'b0000010110001100: out_v[22] = 10'b1011011011;
    16'b0100010100011000: out_v[22] = 10'b1111000111;
    16'b0100110110010100: out_v[22] = 10'b0101011110;
    16'b0100010100001000: out_v[22] = 10'b1000111011;
    16'b0100000110001100: out_v[22] = 10'b0111101000;
    16'b0100010110000100: out_v[22] = 10'b1000110110;
    16'b0100010100010100: out_v[22] = 10'b0100011001;
    16'b0100010100011100: out_v[22] = 10'b0101010100;
    16'b0100000110010100: out_v[22] = 10'b1001001001;
    16'b0100010110010100: out_v[22] = 10'b1001101100;
    16'b0100000100100000: out_v[22] = 10'b0001011011;
    16'b0100010110001100: out_v[22] = 10'b0011011010;
    16'b0100000110000100: out_v[22] = 10'b1100010100;
    16'b0100010110011100: out_v[22] = 10'b0010101100;
    16'b0100000100011000: out_v[22] = 10'b0101010001;
    16'b0000010100010000: out_v[22] = 10'b1111110010;
    16'b0100010100001100: out_v[22] = 10'b1010011010;
    16'b0100000010010100: out_v[22] = 10'b1010001001;
    16'b0000010100001000: out_v[22] = 10'b0011011011;
    16'b0000010100000000: out_v[22] = 10'b1000111010;
    16'b0100000100001000: out_v[22] = 10'b1010001101;
    16'b0000000100000000: out_v[22] = 10'b0111001001;
    16'b0100000110011100: out_v[22] = 10'b0111101110;
    16'b0100010010010100: out_v[22] = 10'b1001110010;
    16'b0000000110000100: out_v[22] = 10'b0001111110;
    16'b0000010100011000: out_v[22] = 10'b0110011000;
    16'b0000100000010100: out_v[22] = 10'b1001101100;
    16'b0100000100010100: out_v[22] = 10'b1101001101;
    16'b0100100000010100: out_v[22] = 10'b1111110011;
    16'b0100000010010000: out_v[22] = 10'b0101011001;
    16'b0000100010010000: out_v[22] = 10'b1001001001;
    16'b0100000000010100: out_v[22] = 10'b1000011110;
    16'b0100010000000000: out_v[22] = 10'b1001001111;
    16'b0100100010010100: out_v[22] = 10'b0111010000;
    16'b0100010110010000: out_v[22] = 10'b1001101010;
    16'b0100010010010000: out_v[22] = 10'b1111011101;
    16'b0100110010010000: out_v[22] = 10'b0100001011;
    16'b0000000000010100: out_v[22] = 10'b0111000011;
    16'b0000000010010000: out_v[22] = 10'b0111010000;
    16'b0000110010010000: out_v[22] = 10'b1100100000;
    16'b0000100010010100: out_v[22] = 10'b1101111000;
    16'b0000010010010000: out_v[22] = 10'b0110110000;
    16'b0100110010010100: out_v[22] = 10'b1110101110;
    16'b0000110010010100: out_v[22] = 10'b1010101001;
    16'b0000100000000000: out_v[22] = 10'b1100101010;
    16'b0100010000011100: out_v[22] = 10'b0110110011;
    16'b0000100010000100: out_v[22] = 10'b0000111000;
    16'b0000110010000100: out_v[22] = 10'b1000101110;
    16'b0100010000011000: out_v[22] = 10'b0011001110;
    16'b0100010010011100: out_v[22] = 10'b1101110010;
    16'b0100010000010010: out_v[22] = 10'b1001010110;
    16'b0100010100010010: out_v[22] = 10'b1110101010;
    16'b0100110000000010: out_v[22] = 10'b1011011111;
    16'b0000010000010010: out_v[22] = 10'b1111100010;
    16'b0100010000000010: out_v[22] = 10'b1011011011;
    16'b0100010100000010: out_v[22] = 10'b0011011100;
    16'b0100110100000010: out_v[22] = 10'b1001110111;
    16'b0000010010000000: out_v[22] = 10'b0110001110;
    16'b0000000010010100: out_v[22] = 10'b0111000101;
    16'b0000010000010100: out_v[22] = 10'b0011100010;
    16'b0100100000011100: out_v[22] = 10'b0110010011;
    16'b0000110000010100: out_v[22] = 10'b1011010110;
    16'b0000000000011000: out_v[22] = 10'b0011010101;
    16'b0100110110011100: out_v[22] = 10'b0111111011;
    16'b0100110010011100: out_v[22] = 10'b0110111011;
    16'b0100110010000100: out_v[22] = 10'b0111101010;
    16'b0100100010000100: out_v[22] = 10'b0100110011;
    16'b0100110100011100: out_v[22] = 10'b0101111011;
    16'b0100110100011000: out_v[22] = 10'b0100110101;
    16'b0100100110001100: out_v[22] = 10'b1001000111;
    16'b0100100100011100: out_v[22] = 10'b1101101100;
    16'b0100100100001100: out_v[22] = 10'b0101101101;
    16'b0100110110000100: out_v[22] = 10'b0100001011;
    16'b0100100010011100: out_v[22] = 10'b0101101110;
    16'b0100100110011100: out_v[22] = 10'b0101011101;
    16'b0100100000001100: out_v[22] = 10'b1110110101;
    16'b0100100000001000: out_v[22] = 10'b1110010011;
    16'b0100010000010100: out_v[22] = 10'b1101100000;
    default: out_v[22] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000000100001: out_v[23] = 10'b1100110011;
    16'b0010100000100100: out_v[23] = 10'b0010001100;
    16'b0010100000000101: out_v[23] = 10'b0001100111;
    16'b0010100000100101: out_v[23] = 10'b1001000000;
    16'b0010000000100001: out_v[23] = 10'b0101001010;
    16'b0000000001100001: out_v[23] = 10'b1101000101;
    16'b0010000000000001: out_v[23] = 10'b0100100001;
    16'b0010100001000001: out_v[23] = 10'b1101010001;
    16'b0000100000100100: out_v[23] = 10'b0001001011;
    16'b0010100000100001: out_v[23] = 10'b1000111001;
    16'b0010000001100001: out_v[23] = 10'b1111010001;
    16'b0010000000100101: out_v[23] = 10'b0110000101;
    16'b0000100000100101: out_v[23] = 10'b0000011010;
    16'b0000000000000001: out_v[23] = 10'b1100001111;
    16'b0010000000000101: out_v[23] = 10'b0010110101;
    16'b0010100001000101: out_v[23] = 10'b0101110011;
    16'b0010100001100001: out_v[23] = 10'b1111111010;
    16'b0000100001100101: out_v[23] = 10'b1000011110;
    16'b0010000000101001: out_v[23] = 10'b0101010011;
    16'b0000000000100101: out_v[23] = 10'b0001100100;
    16'b0010000000000000: out_v[23] = 10'b1111100100;
    16'b0000100001000100: out_v[23] = 10'b0001001111;
    16'b0000000000100000: out_v[23] = 10'b1000101110;
    16'b0000100001100100: out_v[23] = 10'b1010101101;
    16'b0000100000000100: out_v[23] = 10'b0111010001;
    16'b0010100001100101: out_v[23] = 10'b0100101001;
    16'b0010000000100000: out_v[23] = 10'b0101100011;
    16'b0000000000000000: out_v[23] = 10'b0010001111;
    16'b0010000001000001: out_v[23] = 10'b0000010111;
    16'b0010000001100101: out_v[23] = 10'b1101110111;
    16'b0010100000000001: out_v[23] = 10'b1100110001;
    16'b0000000001100000: out_v[23] = 10'b0011111001;
    16'b0000000000100100: out_v[23] = 10'b0111110100;
    16'b0000000001100101: out_v[23] = 10'b1110000100;
    16'b0000000001100100: out_v[23] = 10'b1011100110;
    16'b0000000001000000: out_v[23] = 10'b0010110110;
    16'b0000000000000100: out_v[23] = 10'b1000101010;
    16'b0000000001000001: out_v[23] = 10'b1010110111;
    16'b0000100001101100: out_v[23] = 10'b1101010011;
    16'b0000100000101000: out_v[23] = 10'b1110010100;
    16'b0000000001101000: out_v[23] = 10'b1000011100;
    16'b0000100001000000: out_v[23] = 10'b0001011111;
    16'b0000000000110000: out_v[23] = 10'b0000110100;
    16'b0000000001010000: out_v[23] = 10'b1010010100;
    16'b0000100001100000: out_v[23] = 10'b1010100110;
    16'b0000100001101000: out_v[23] = 10'b0011010111;
    16'b0000000000010000: out_v[23] = 10'b1111000101;
    16'b0000100001100001: out_v[23] = 10'b0000111111;
    16'b0000000001000100: out_v[23] = 10'b1111010100;
    16'b0000100001111000: out_v[23] = 10'b1111101011;
    16'b0000000000101000: out_v[23] = 10'b1010011100;
    16'b0000000001101100: out_v[23] = 10'b0011010011;
    16'b0000000001001000: out_v[23] = 10'b0110110000;
    16'b0000100000101100: out_v[23] = 10'b1011101100;
    16'b0000001001000000: out_v[23] = 10'b0111100110;
    16'b0000100000100000: out_v[23] = 10'b1111001100;
    16'b0000000000101100: out_v[23] = 10'b1111101101;
    16'b0000100001110100: out_v[23] = 10'b0011110111;
    16'b0000001000000000: out_v[23] = 10'b0000001011;
    16'b0000101000100100: out_v[23] = 10'b1111110011;
    16'b0000000100100000: out_v[23] = 10'b1011011011;
    16'b0010100001100100: out_v[23] = 10'b0001001110;
    16'b0000000101100000: out_v[23] = 10'b1111111111;
    16'b0000100101100100: out_v[23] = 10'b0001111011;
    16'b0010000001000000: out_v[23] = 10'b1101010000;
    16'b0010000001000010: out_v[23] = 10'b0101110110;
    16'b0010000001000011: out_v[23] = 10'b1000101001;
    16'b0010000001100000: out_v[23] = 10'b0100010000;
    16'b0000100001000001: out_v[23] = 10'b0010101100;
    16'b0000100001000101: out_v[23] = 10'b1001101110;
    16'b0000000001000101: out_v[23] = 10'b1111100111;
    16'b0000100000000101: out_v[23] = 10'b1001111111;
    16'b0010000001000101: out_v[23] = 10'b0110010010;
    16'b0000100000000000: out_v[23] = 10'b1111001010;
    16'b0000100000100001: out_v[23] = 10'b0111100110;
    16'b0010000000001001: out_v[23] = 10'b0011100100;
    16'b0000000001101001: out_v[23] = 10'b0110111110;
    16'b0010000001001001: out_v[23] = 10'b1011010010;
    16'b0000000000001000: out_v[23] = 10'b1001100011;
    16'b0000000000001001: out_v[23] = 10'b1111110011;
    16'b0010000001101001: out_v[23] = 10'b1011001110;
    16'b0000000001001001: out_v[23] = 10'b1111101010;
    16'b0000000000101001: out_v[23] = 10'b1110111011;
    16'b0010000000001000: out_v[23] = 10'b1011100001;
    16'b0000000001000011: out_v[23] = 10'b0111100011;
    16'b0000001001000011: out_v[23] = 10'b1010011011;
    16'b0010000000000011: out_v[23] = 10'b1110100110;
    16'b0000001001000001: out_v[23] = 10'b1011110100;
    16'b0000000001000010: out_v[23] = 10'b1010100100;
    16'b0000000000000011: out_v[23] = 10'b0001110110;
    16'b0000000000000101: out_v[23] = 10'b0101011010;
    16'b0010000000000010: out_v[23] = 10'b1000101011;
    default: out_v[23] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1011000000000000: out_v[24] = 10'b0100001001;
    16'b0011000000000001: out_v[24] = 10'b1101011010;
    16'b1001000000000001: out_v[24] = 10'b0111110010;
    16'b1001100000000000: out_v[24] = 10'b0000000101;
    16'b1010000000000000: out_v[24] = 10'b0011000101;
    16'b1001000000000000: out_v[24] = 10'b0010111001;
    16'b1000000000000000: out_v[24] = 10'b0010100011;
    16'b0010000000000000: out_v[24] = 10'b0010001001;
    16'b0011000000000000: out_v[24] = 10'b0000001101;
    16'b0011000001000000: out_v[24] = 10'b1001010010;
    16'b0001000000000000: out_v[24] = 10'b0010011010;
    16'b1011000000000001: out_v[24] = 10'b0000100001;
    16'b0010000000000001: out_v[24] = 10'b0010001011;
    16'b1011100000000000: out_v[24] = 10'b1100000001;
    16'b1000100000000001: out_v[24] = 10'b0001010011;
    16'b0000000000000000: out_v[24] = 10'b0011101011;
    16'b1000000000000001: out_v[24] = 10'b1001100001;
    16'b1001100000000001: out_v[24] = 10'b1010010111;
    16'b1011100000000001: out_v[24] = 10'b1001110011;
    16'b0001100000000000: out_v[24] = 10'b1101011011;
    16'b1000100000000000: out_v[24] = 10'b1100001101;
    16'b1001100000001000: out_v[24] = 10'b0111101001;
    16'b0001000000000001: out_v[24] = 10'b0101011111;
    16'b0010000001000000: out_v[24] = 10'b0111000111;
    16'b1011000001000000: out_v[24] = 10'b0000111101;
    16'b0010000101000000: out_v[24] = 10'b0010010101;
    16'b1011100100000000: out_v[24] = 10'b1101011010;
    16'b1011000101000000: out_v[24] = 10'b0111010111;
    16'b0000000101000000: out_v[24] = 10'b0011010011;
    16'b0000000101000001: out_v[24] = 10'b1001110010;
    16'b0000000100000000: out_v[24] = 10'b1100100100;
    16'b0000000100000001: out_v[24] = 10'b1110100000;
    16'b0001000101000000: out_v[24] = 10'b1000110100;
    16'b0001000100000000: out_v[24] = 10'b0101010110;
    16'b0011000101000000: out_v[24] = 10'b1000110011;
    16'b0000000001000000: out_v[24] = 10'b0101011001;
    16'b1000000101000000: out_v[24] = 10'b0110110000;
    16'b1001000101000000: out_v[24] = 10'b0101000110;
    16'b1011000100000000: out_v[24] = 10'b1101100011;
    16'b0010000100000000: out_v[24] = 10'b0101001010;
    16'b0001000001000000: out_v[24] = 10'b1000011001;
    16'b0011100101000000: out_v[24] = 10'b1011101100;
    16'b0001100101000000: out_v[24] = 10'b0011000110;
    16'b0011000100000000: out_v[24] = 10'b0100111100;
    16'b1001000100000000: out_v[24] = 10'b0101011011;
    16'b1000000100000000: out_v[24] = 10'b1011010100;
    16'b1010000100000000: out_v[24] = 10'b1101100111;
    16'b0010100101000000: out_v[24] = 10'b0110101110;
    16'b1010000101000000: out_v[24] = 10'b0111001010;
    16'b0001010101000000: out_v[24] = 10'b1100101101;
    16'b0000010101000000: out_v[24] = 10'b0111000110;
    16'b0000000001000001: out_v[24] = 10'b0100101101;
    16'b0001000001000001: out_v[24] = 10'b1101000101;
    16'b0011000001000001: out_v[24] = 10'b0000100111;
    16'b0010000001000001: out_v[24] = 10'b0011111011;
    16'b0011100000000000: out_v[24] = 10'b0010001110;
    16'b1000000001000001: out_v[24] = 10'b0011100110;
    16'b0000000000000001: out_v[24] = 10'b1001111111;
    16'b0001000101000001: out_v[24] = 10'b1011011010;
    16'b1000000101000001: out_v[24] = 10'b1100101000;
    16'b1001000001000001: out_v[24] = 10'b0111011111;
    16'b1011000001000001: out_v[24] = 10'b1000001110;
    16'b0010000101000001: out_v[24] = 10'b0010001110;
    16'b1010000001000000: out_v[24] = 10'b0100110010;
    16'b1010000101000001: out_v[24] = 10'b1101001010;
    16'b1000000001000000: out_v[24] = 10'b1001101000;
    16'b1010100001000000: out_v[24] = 10'b1110010010;
    16'b1010100101000000: out_v[24] = 10'b0111100000;
    16'b1011100101000000: out_v[24] = 10'b1011010011;
    16'b1000000111000000: out_v[24] = 10'b1101001101;
    16'b1010000011000000: out_v[24] = 10'b1000011110;
    16'b1010000111000000: out_v[24] = 10'b0101011111;
    16'b1001000001000000: out_v[24] = 10'b0110100011;
    16'b1001000101000001: out_v[24] = 10'b1011111011;
    16'b1010000000000001: out_v[24] = 10'b1111000110;
    16'b1000000111000001: out_v[24] = 10'b0100110000;
    16'b1010000100001001: out_v[24] = 10'b0011000110;
    16'b1011000010001000: out_v[24] = 10'b1011010101;
    16'b1010000010000001: out_v[24] = 10'b0110101101;
    16'b1000000100000001: out_v[24] = 10'b0110111111;
    16'b1000000010000000: out_v[24] = 10'b0010110100;
    16'b0000000010000000: out_v[24] = 10'b0111111001;
    16'b1010000010000000: out_v[24] = 10'b0111011011;
    16'b1010000100000001: out_v[24] = 10'b0110111000;
    16'b1010000000001001: out_v[24] = 10'b0011110011;
    16'b1000000010001000: out_v[24] = 10'b1101011111;
    16'b1000000110000000: out_v[24] = 10'b0011100010;
    16'b1011000000001000: out_v[24] = 10'b0101011111;
    16'b0000000110000001: out_v[24] = 10'b0000110111;
    16'b0010000100000001: out_v[24] = 10'b1010011100;
    16'b1010000010001000: out_v[24] = 10'b0100100110;
    16'b1010000000001000: out_v[24] = 10'b1101110110;
    16'b0010000010000000: out_v[24] = 10'b1111101010;
    16'b1011000000001010: out_v[24] = 10'b0001110101;
    16'b0000000110000000: out_v[24] = 10'b1000101010;
    16'b1010000110000001: out_v[24] = 10'b0110110101;
    16'b1000000110000001: out_v[24] = 10'b0111011101;
    16'b1010000010001001: out_v[24] = 10'b1111011111;
    16'b1000000000001000: out_v[24] = 10'b0011001101;
    16'b1010000111000001: out_v[24] = 10'b1100111110;
    16'b1011000101000001: out_v[24] = 10'b1101010000;
    16'b1010000001000001: out_v[24] = 10'b1101110011;
    16'b1000000101000010: out_v[24] = 10'b1101000111;
    16'b1010000110000000: out_v[24] = 10'b1000001010;
    16'b1000000011000000: out_v[24] = 10'b1001101011;
    16'b0000000011000000: out_v[24] = 10'b1101001101;
    16'b1011000100000010: out_v[24] = 10'b1001101110;
    16'b0000000111000000: out_v[24] = 10'b1101100101;
    16'b1010000011000001: out_v[24] = 10'b1110010011;
    16'b1011000001000010: out_v[24] = 10'b1001001110;
    16'b1000000001000010: out_v[24] = 10'b1001100001;
    16'b1011000101000010: out_v[24] = 10'b1001010111;
    16'b1011000101100010: out_v[24] = 10'b1101111110;
    default: out_v[24] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1001000000000001: out_v[25] = 10'b1101001100;
    16'b1100010100000001: out_v[25] = 10'b0111111010;
    16'b1100010100001001: out_v[25] = 10'b1111010011;
    16'b1101000000001001: out_v[25] = 10'b1011000011;
    16'b1101000100001000: out_v[25] = 10'b1000000001;
    16'b1100010100000000: out_v[25] = 10'b0100111111;
    16'b1100010000001001: out_v[25] = 10'b0100111000;
    16'b1000010100000000: out_v[25] = 10'b0111110011;
    16'b1100010000000001: out_v[25] = 10'b1000101011;
    16'b1101000000000001: out_v[25] = 10'b0001100001;
    16'b1101000100001001: out_v[25] = 10'b1000100011;
    16'b1100000000000001: out_v[25] = 10'b0000100001;
    16'b1101000100000000: out_v[25] = 10'b1001100001;
    16'b1101010000001001: out_v[25] = 10'b0011001101;
    16'b1101010000000001: out_v[25] = 10'b1011000101;
    16'b1101010100000001: out_v[25] = 10'b1010001000;
    16'b1100010100001000: out_v[25] = 10'b0101010000;
    16'b1100010000000000: out_v[25] = 10'b0010011101;
    16'b0100010000000001: out_v[25] = 10'b0000101010;
    16'b0101000100001000: out_v[25] = 10'b0011100111;
    16'b0100010100000000: out_v[25] = 10'b0101001111;
    16'b0000010000000001: out_v[25] = 10'b0010000111;
    16'b1101010100001001: out_v[25] = 10'b1000000011;
    16'b1101000100000001: out_v[25] = 10'b0110011111;
    16'b1000010000000001: out_v[25] = 10'b0010111101;
    16'b1100000000001001: out_v[25] = 10'b1111010011;
    16'b0001000000000001: out_v[25] = 10'b1010001010;
    16'b1101010100001000: out_v[25] = 10'b0001001001;
    16'b0101010100000000: out_v[25] = 10'b1000000110;
    16'b1101010100000000: out_v[25] = 10'b1000010011;
    16'b1100010000001000: out_v[25] = 10'b1011010010;
    16'b0101000100000000: out_v[25] = 10'b1001001101;
    16'b0100000000000001: out_v[25] = 10'b0100101011;
    16'b1000010000000000: out_v[25] = 10'b1011000110;
    16'b1101110100001000: out_v[25] = 10'b1001001011;
    16'b1000010000001001: out_v[25] = 10'b0111111010;
    16'b0000000100001000: out_v[25] = 10'b0101000101;
    16'b0000000100000000: out_v[25] = 10'b1100011100;
    16'b0000000100000001: out_v[25] = 10'b1010110111;
    16'b0000000000001000: out_v[25] = 10'b0011100011;
    16'b0000000000000000: out_v[25] = 10'b0011110011;
    16'b0000000100001001: out_v[25] = 10'b1010010011;
    16'b1000000100000001: out_v[25] = 10'b0110001000;
    16'b1000000100000000: out_v[25] = 10'b0100101110;
    16'b0000100000000000: out_v[25] = 10'b0000111010;
    16'b0000000000000001: out_v[25] = 10'b0000001100;
    16'b0001000100000000: out_v[25] = 10'b0110001001;
    16'b0100000100001000: out_v[25] = 10'b1011100100;
    16'b0101010100001000: out_v[25] = 10'b0010010110;
    16'b0101010000000000: out_v[25] = 10'b0101010110;
    16'b0000000000001001: out_v[25] = 10'b1110011100;
    16'b1100000100001000: out_v[25] = 10'b0111001110;
    16'b1001000100001000: out_v[25] = 10'b1101111110;
    16'b0001000100001000: out_v[25] = 10'b1000101000;
    16'b0100010100001000: out_v[25] = 10'b1100100100;
    16'b0100000100000000: out_v[25] = 10'b1111100110;
    16'b0001000100000001: out_v[25] = 10'b1100110100;
    16'b0100010000000000: out_v[25] = 10'b1111100111;
    16'b1001000100000000: out_v[25] = 10'b0001001100;
    16'b1000000100001000: out_v[25] = 10'b1111001110;
    16'b0100000000001000: out_v[25] = 10'b1000111111;
    16'b1100000100000000: out_v[25] = 10'b1001110110;
    16'b1000000000000000: out_v[25] = 10'b0010101010;
    16'b1100000000000000: out_v[25] = 10'b1001011100;
    16'b0100010000001000: out_v[25] = 10'b1100100101;
    16'b0100000000000000: out_v[25] = 10'b1111110100;
    16'b0100000100000001: out_v[25] = 10'b0100011011;
    16'b1001000000001001: out_v[25] = 10'b1110100010;
    16'b0001000000000000: out_v[25] = 10'b0111011110;
    16'b1000000000000001: out_v[25] = 10'b1101100000;
    16'b0101000000000001: out_v[25] = 10'b1100010101;
    16'b0101010000000001: out_v[25] = 10'b1101011010;
    16'b0001000000001001: out_v[25] = 10'b1010001011;
    16'b1001000100000001: out_v[25] = 10'b0110001111;
    16'b0001000100001001: out_v[25] = 10'b0011001010;
    16'b0001000000001000: out_v[25] = 10'b1111110000;
    16'b1101000000000000: out_v[25] = 10'b0010110011;
    16'b0101000000000000: out_v[25] = 10'b1010010011;
    16'b1101110100000000: out_v[25] = 10'b1011100111;
    16'b1100000100000001: out_v[25] = 10'b1111100000;
    16'b1101010000000000: out_v[25] = 10'b0000111010;
    16'b1101110100000001: out_v[25] = 10'b1011110111;
    16'b1100110100000000: out_v[25] = 10'b1111010001;
    16'b0101000100000001: out_v[25] = 10'b1101100100;
    16'b0101010000001000: out_v[25] = 10'b1110111011;
    16'b0111010000000000: out_v[25] = 10'b1100010010;
    16'b1101010000001000: out_v[25] = 10'b0001011000;
    16'b1100100100000000: out_v[25] = 10'b1001111111;
    16'b0101010100000001: out_v[25] = 10'b0010010100;
    16'b1001000000000000: out_v[25] = 10'b1110110000;
    16'b1001100000000001: out_v[25] = 10'b1111011011;
    16'b1000100100000001: out_v[25] = 10'b1111001010;
    16'b1000100100000000: out_v[25] = 10'b0100100100;
    16'b1000100000000001: out_v[25] = 10'b1000100111;
    16'b1100100000000001: out_v[25] = 10'b0011100100;
    16'b1000000000001001: out_v[25] = 10'b0000100100;
    16'b1100100100000001: out_v[25] = 10'b1110110110;
    16'b0000100100000000: out_v[25] = 10'b1011110100;
    16'b0000100000000001: out_v[25] = 10'b1010111010;
    16'b1000100000001001: out_v[25] = 10'b1001111110;
    16'b1100110000000001: out_v[25] = 10'b1111101011;
    16'b1100000000001000: out_v[25] = 10'b1101100011;
    16'b1101000000001000: out_v[25] = 10'b1111011000;
    16'b0000010100000000: out_v[25] = 10'b0101110011;
    16'b1001010100000001: out_v[25] = 10'b1100001000;
    16'b1001010000000000: out_v[25] = 10'b1111000010;
    16'b1000000100001001: out_v[25] = 10'b0110011000;
    16'b1111010000000000: out_v[25] = 10'b1011001011;
    default: out_v[25] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001000000001000: out_v[26] = 10'b1111010000;
    16'b1000000000001010: out_v[26] = 10'b0110001000;
    16'b1001000001001010: out_v[26] = 10'b0001001010;
    16'b0001000000000010: out_v[26] = 10'b0011011001;
    16'b1001000001111010: out_v[26] = 10'b1111011011;
    16'b1000000000000010: out_v[26] = 10'b0110001011;
    16'b1001000001000010: out_v[26] = 10'b1000110111;
    16'b1000000001000010: out_v[26] = 10'b1101011001;
    16'b0001000001110010: out_v[26] = 10'b1011001110;
    16'b1001000000001010: out_v[26] = 10'b1000100101;
    16'b1000000001011010: out_v[26] = 10'b1000011100;
    16'b1000000001000011: out_v[26] = 10'b0110011111;
    16'b0001000001000010: out_v[26] = 10'b1111000111;
    16'b0001000001000000: out_v[26] = 10'b0011001101;
    16'b0001000001001010: out_v[26] = 10'b1111100011;
    16'b1001000000000010: out_v[26] = 10'b0111011110;
    16'b1001000001010010: out_v[26] = 10'b0000110001;
    16'b1001000001110010: out_v[26] = 10'b0100111001;
    16'b1000000001010010: out_v[26] = 10'b1100110110;
    16'b1000000001001010: out_v[26] = 10'b0010011000;
    16'b0001100001110010: out_v[26] = 10'b1011110011;
    16'b0001000001110000: out_v[26] = 10'b1010011001;
    16'b0001000000001010: out_v[26] = 10'b0010110101;
    16'b1000000000000011: out_v[26] = 10'b1010110011;
    16'b1001100001110010: out_v[26] = 10'b1100100101;
    16'b0001000001111010: out_v[26] = 10'b1001011110;
    16'b0001000001010010: out_v[26] = 10'b0010111011;
    16'b0001000000000000: out_v[26] = 10'b1010100011;
    16'b1001000001010011: out_v[26] = 10'b1001011110;
    16'b0001000001001000: out_v[26] = 10'b0111110111;
    16'b1001100001111010: out_v[26] = 10'b0000001011;
    16'b1100000000000010: out_v[26] = 10'b1010111001;
    16'b1001000001000011: out_v[26] = 10'b0111111110;
    16'b1001000001011010: out_v[26] = 10'b0010100011;
    16'b0001000001010000: out_v[26] = 10'b1000101011;
    16'b1100000000001010: out_v[26] = 10'b1001111011;
    16'b0100000000001000: out_v[26] = 10'b1011001010;
    16'b1101000000000010: out_v[26] = 10'b1001101010;
    16'b0000000000000000: out_v[26] = 10'b1011000011;
    16'b1101000000000000: out_v[26] = 10'b0011010010;
    16'b1100000000000000: out_v[26] = 10'b1101110000;
    16'b0000000000001000: out_v[26] = 10'b1011000011;
    16'b0000000000000010: out_v[26] = 10'b0010010011;
    16'b0100000000000010: out_v[26] = 10'b0100011010;
    16'b0100000000000000: out_v[26] = 10'b1001100101;
    16'b0100000000001010: out_v[26] = 10'b1000011010;
    16'b0101000000000000: out_v[26] = 10'b0110011100;
    16'b0000000000001010: out_v[26] = 10'b0111100101;
    16'b1101100000101010: out_v[26] = 10'b1110100111;
    16'b0100000001011000: out_v[26] = 10'b0011100101;
    16'b1001100001101010: out_v[26] = 10'b1100100100;
    16'b1100000001101010: out_v[26] = 10'b1000111111;
    16'b1101100000001010: out_v[26] = 10'b1111110110;
    16'b1100000001100010: out_v[26] = 10'b1100000011;
    16'b1100000001001010: out_v[26] = 10'b1010110110;
    16'b1100100000001010: out_v[26] = 10'b0010100001;
    16'b0100000001111000: out_v[26] = 10'b1010001011;
    16'b0100000001100000: out_v[26] = 10'b0101101101;
    16'b1100000000001000: out_v[26] = 10'b1101100011;
    16'b0100000001010000: out_v[26] = 10'b0100000100;
    16'b0101000000001000: out_v[26] = 10'b1101001000;
    16'b1100100001101010: out_v[26] = 10'b0000000111;
    16'b1001100000001010: out_v[26] = 10'b1001010111;
    16'b1100000000101000: out_v[26] = 10'b0100001101;
    16'b0100000000101000: out_v[26] = 10'b0011011111;
    16'b1100000001111010: out_v[26] = 10'b1010111110;
    16'b1100000000101010: out_v[26] = 10'b1000101110;
    16'b0100000001101000: out_v[26] = 10'b0000111110;
    16'b1100100001111010: out_v[26] = 10'b0110110101;
    16'b1101000000101010: out_v[26] = 10'b1010010110;
    16'b1100000001101000: out_v[26] = 10'b1110100011;
    16'b1001100000100010: out_v[26] = 10'b0001011110;
    16'b1001100000101010: out_v[26] = 10'b0000110110;
    16'b0100000001001000: out_v[26] = 10'b0010100100;
    16'b1101000000001000: out_v[26] = 10'b0010011100;
    16'b1101000000001010: out_v[26] = 10'b1111111100;
    16'b1100100001011010: out_v[26] = 10'b0111011010;
    16'b0101000000001010: out_v[26] = 10'b0110100000;
    16'b1100000001000010: out_v[26] = 10'b1010110011;
    16'b1100100000101010: out_v[26] = 10'b1101011011;
    16'b1100000001001000: out_v[26] = 10'b0011100101;
    16'b1101100001101010: out_v[26] = 10'b0010111000;
    16'b1100000001011010: out_v[26] = 10'b1011011110;
    16'b0100000000011000: out_v[26] = 10'b1110100111;
    16'b0001100001000000: out_v[26] = 10'b1111001101;
    16'b1001100001001010: out_v[26] = 10'b0110111011;
    16'b0101100000001000: out_v[26] = 10'b0010101111;
    16'b0001100000000000: out_v[26] = 10'b0000011110;
    16'b0101100000000000: out_v[26] = 10'b1011001111;
    16'b0001100001100000: out_v[26] = 10'b1010001101;
    16'b0001100001000010: out_v[26] = 10'b0011011011;
    16'b0001100000001000: out_v[26] = 10'b1001000100;
    16'b0001100000000010: out_v[26] = 10'b1110000010;
    16'b0101000000000010: out_v[26] = 10'b1101011000;
    16'b0001100001111010: out_v[26] = 10'b0110110010;
    16'b0001100000001010: out_v[26] = 10'b0001001110;
    16'b0101100000001010: out_v[26] = 10'b0101110010;
    16'b1101100001001010: out_v[26] = 10'b1000101111;
    16'b0001100001001000: out_v[26] = 10'b0110100010;
    16'b0001100001001010: out_v[26] = 10'b0011101010;
    16'b0001100001101010: out_v[26] = 10'b0110110011;
    16'b1101100000000010: out_v[26] = 10'b1101000100;
    16'b1001100001000010: out_v[26] = 10'b0111001001;
    16'b1001100000000010: out_v[26] = 10'b1000110100;
    16'b0001100001100010: out_v[26] = 10'b1010110111;
    16'b1100000000001011: out_v[26] = 10'b1111110110;
    16'b0100000000001001: out_v[26] = 10'b0110011110;
    16'b1101100000001000: out_v[26] = 10'b1001100111;
    16'b1001000000001000: out_v[26] = 10'b1101000100;
    16'b0100100000001000: out_v[26] = 10'b0100111010;
    16'b1100000000011010: out_v[26] = 10'b1011110010;
    16'b1100000000000011: out_v[26] = 10'b0100110001;
    16'b0000100000001000: out_v[26] = 10'b0001010101;
    16'b0101000000000001: out_v[26] = 10'b1010110110;
    16'b1001000000000011: out_v[26] = 10'b0001110110;
    16'b1101000000000011: out_v[26] = 10'b1000111011;
    16'b0101000000000011: out_v[26] = 10'b1000100010;
    16'b1000000000001011: out_v[26] = 10'b0100111010;
    16'b1000000000000001: out_v[26] = 10'b0110001111;
    16'b1100000000000001: out_v[26] = 10'b1111101011;
    16'b0000000000001001: out_v[26] = 10'b1000100000;
    16'b0001000000000001: out_v[26] = 10'b0001110110;
    16'b1101000001000010: out_v[26] = 10'b1011101000;
    16'b1101000001001010: out_v[26] = 10'b1111010001;
    16'b1100000001010010: out_v[26] = 10'b1110011110;
    16'b1100000001000000: out_v[26] = 10'b0001001011;
    16'b1100000001110010: out_v[26] = 10'b1000110010;
    16'b1000000000000000: out_v[26] = 10'b0111111100;
    16'b1101000000001011: out_v[26] = 10'b0110011100;
    16'b0101000001001010: out_v[26] = 10'b0100011111;
    16'b0101000000001001: out_v[26] = 10'b0111010111;
    16'b1000000000001000: out_v[26] = 10'b1000101110;
    default: out_v[26] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100000000000000: out_v[27] = 10'b0100010111;
    16'b1100000000000001: out_v[27] = 10'b0100010111;
    16'b0000000000000001: out_v[27] = 10'b1111010000;
    16'b0000000000000101: out_v[27] = 10'b1000110111;
    16'b0100000000000001: out_v[27] = 10'b0101010001;
    16'b0000000000000000: out_v[27] = 10'b0000011110;
    16'b0100000000000101: out_v[27] = 10'b1111110010;
    16'b1000000000000101: out_v[27] = 10'b0000011101;
    16'b0000000000000100: out_v[27] = 10'b0100110010;
    16'b1000000000000001: out_v[27] = 10'b0110110101;
    16'b1100000000000100: out_v[27] = 10'b0101010100;
    16'b0100000000000100: out_v[27] = 10'b0001110010;
    16'b1100000000000101: out_v[27] = 10'b0100101011;
    16'b1100000000000000: out_v[27] = 10'b0100110010;
    16'b1000000000000000: out_v[27] = 10'b0110110000;
    16'b0100000000100000: out_v[27] = 10'b1001010100;
    16'b1000000000000100: out_v[27] = 10'b1010001000;
    16'b0000000000001000: out_v[27] = 10'b1110011001;
    16'b0000000000010000: out_v[27] = 10'b1100000100;
    16'b0100000000010000: out_v[27] = 10'b1010101000;
    16'b0100000000100001: out_v[27] = 10'b1001001100;
    16'b0000000000100000: out_v[27] = 10'b0101000011;
    16'b0000000000100001: out_v[27] = 10'b1101110000;
    16'b0000000000000010: out_v[27] = 10'b1011000010;
    16'b0000000010000000: out_v[27] = 10'b1000001000;
    16'b0000000000010010: out_v[27] = 10'b1110001000;
    16'b0100000000000010: out_v[27] = 10'b1010001011;
    16'b0001000000000000: out_v[27] = 10'b0110010100;
    default: out_v[27] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000001000001000: out_v[28] = 10'b0001011101;
    16'b0000000010111000: out_v[28] = 10'b0100000111;
    16'b0000100010101000: out_v[28] = 10'b1101001110;
    16'b0000000000101000: out_v[28] = 10'b1001011010;
    16'b0000000010001000: out_v[28] = 10'b1110110010;
    16'b0000000000001000: out_v[28] = 10'b0011101001;
    16'b0000000010101000: out_v[28] = 10'b0000101100;
    16'b0000000000000000: out_v[28] = 10'b0100101100;
    16'b0000001010001000: out_v[28] = 10'b0011001010;
    16'b0000001000101000: out_v[28] = 10'b0101100111;
    16'b0000001010101000: out_v[28] = 10'b1101000100;
    16'b0000000010000000: out_v[28] = 10'b1011000001;
    16'b0000100000101000: out_v[28] = 10'b0000110001;
    16'b0000100000100000: out_v[28] = 10'b1110100001;
    16'b0000000000100000: out_v[28] = 10'b0010101011;
    16'b0000100000001000: out_v[28] = 10'b1011111101;
    16'b0000001010111000: out_v[28] = 10'b1111101100;
    16'b0000000010100000: out_v[28] = 10'b0100101101;
    16'b0000000000111000: out_v[28] = 10'b0000001101;
    16'b0000100000000000: out_v[28] = 10'b1110100010;
    16'b0000001000000000: out_v[28] = 10'b0100110111;
    16'b0000001010000000: out_v[28] = 10'b1001010011;
    16'b0000001010100000: out_v[28] = 10'b0100010101;
    16'b0000000000110000: out_v[28] = 10'b1101010101;
    16'b0000001000100000: out_v[28] = 10'b0110000000;
    16'b0000100010001000: out_v[28] = 10'b1111000110;
    16'b0000000010110000: out_v[28] = 10'b1000111011;
    16'b0000000010011000: out_v[28] = 10'b1011011011;
    16'b0000001000111000: out_v[28] = 10'b0001001011;
    16'b0000101010001000: out_v[28] = 10'b1111100001;
    16'b0000101010000000: out_v[28] = 10'b1110010010;
    16'b0000101000000000: out_v[28] = 10'b1100011011;
    16'b0000000100010000: out_v[28] = 10'b0001001011;
    16'b0000010010000000: out_v[28] = 10'b0011100111;
    16'b0000010010001000: out_v[28] = 10'b0101111110;
    16'b0000010000000000: out_v[28] = 10'b1010101001;
    16'b0000100010000000: out_v[28] = 10'b0110100101;
    16'b0000000100000000: out_v[28] = 10'b0010110000;
    16'b0000110010000000: out_v[28] = 10'b0101111011;
    16'b0000000110010000: out_v[28] = 10'b1110000110;
    16'b0000000110000000: out_v[28] = 10'b1111000101;
    16'b0000000100110000: out_v[28] = 10'b1011000101;
    16'b0000000110110000: out_v[28] = 10'b1011000010;
    16'b0000110010001000: out_v[28] = 10'b0111001000;
    16'b0000100110010000: out_v[28] = 10'b0001111011;
    16'b0000001100110000: out_v[28] = 10'b1001010110;
    16'b0000001000110000: out_v[28] = 10'b1110001010;
    16'b0000001010110000: out_v[28] = 10'b1001111111;
    16'b0000001110000000: out_v[28] = 10'b1001110111;
    16'b0000011010000000: out_v[28] = 10'b1001100101;
    16'b0000101000001000: out_v[28] = 10'b0100101011;
    default: out_v[28] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1000010100100001: out_v[29] = 10'b0101011101;
    16'b1010010100000001: out_v[29] = 10'b1001000011;
    16'b0010010100000001: out_v[29] = 10'b1100100010;
    16'b1010010000000000: out_v[29] = 10'b0100011000;
    16'b0010010100100001: out_v[29] = 10'b0111011111;
    16'b0000010100100001: out_v[29] = 10'b0110000111;
    16'b1010000110000001: out_v[29] = 10'b1011100110;
    16'b0000010000000000: out_v[29] = 10'b1100101011;
    16'b1010000000000000: out_v[29] = 10'b0100001101;
    16'b1010010110000001: out_v[29] = 10'b0101100110;
    16'b1010010100100001: out_v[29] = 10'b1010100101;
    16'b1000010000000000: out_v[29] = 10'b0010011111;
    16'b1010010100000000: out_v[29] = 10'b0100100010;
    16'b0010010100000000: out_v[29] = 10'b1110000111;
    16'b0000010100100000: out_v[29] = 10'b0010110101;
    16'b1010000100000001: out_v[29] = 10'b1110100011;
    16'b0010010000000000: out_v[29] = 10'b0100001011;
    16'b1010010000000001: out_v[29] = 10'b0011010101;
    16'b1000010000100000: out_v[29] = 10'b0111010010;
    16'b1010000100000000: out_v[29] = 10'b1110000110;
    16'b1010010110100001: out_v[29] = 10'b1011100111;
    16'b1000010100000001: out_v[29] = 10'b1010100100;
    16'b0010010000000001: out_v[29] = 10'b1100100001;
    16'b1000010100100000: out_v[29] = 10'b1000101111;
    16'b1010010000100000: out_v[29] = 10'b0000111111;
    16'b1000000000000000: out_v[29] = 10'b1100001100;
    16'b0010010000100000: out_v[29] = 10'b1100010011;
    16'b1010010010000001: out_v[29] = 10'b1001010100;
    16'b0000010000100000: out_v[29] = 10'b1001000100;
    16'b1010010100100000: out_v[29] = 10'b1010010101;
    16'b0010000000000000: out_v[29] = 10'b0101100100;
    16'b1010010010100000: out_v[29] = 10'b0001111110;
    16'b0000000000000000: out_v[29] = 10'b0001010001;
    16'b0000000000000001: out_v[29] = 10'b0010011011;
    16'b0010010010100000: out_v[29] = 10'b1011011010;
    16'b0010000010100000: out_v[29] = 10'b1010001111;
    16'b0000000100000001: out_v[29] = 10'b0010011111;
    16'b0000010000000001: out_v[29] = 10'b1101011110;
    16'b1000010010100000: out_v[29] = 10'b1011101110;
    16'b0010000000100000: out_v[29] = 10'b0001010110;
    16'b0000010010100000: out_v[29] = 10'b0101000000;
    16'b0000010100000001: out_v[29] = 10'b0010101110;
    16'b1010000000100000: out_v[29] = 10'b0010010101;
    16'b1010000010000000: out_v[29] = 10'b0001011110;
    16'b0000000000100000: out_v[29] = 10'b1001100100;
    16'b1000000000100000: out_v[29] = 10'b1100000000;
    16'b0010000010000000: out_v[29] = 10'b0000101101;
    16'b1010000010100000: out_v[29] = 10'b0000101101;
    16'b1001010000000000: out_v[29] = 10'b0000011010;
    16'b1010010010000000: out_v[29] = 10'b0101101101;
    16'b0010000100000001: out_v[29] = 10'b0101100000;
    16'b0000010100000000: out_v[29] = 10'b1101100000;
    16'b0000000100000000: out_v[29] = 10'b0000011001;
    16'b0000000100100001: out_v[29] = 10'b0111011110;
    16'b1000010100000000: out_v[29] = 10'b1001011100;
    16'b0000000110000001: out_v[29] = 10'b1010101011;
    16'b0000000110000000: out_v[29] = 10'b1010101001;
    16'b0000000010000000: out_v[29] = 10'b1110010101;
    16'b1000010000000001: out_v[29] = 10'b1100011100;
    16'b0010000100100001: out_v[29] = 10'b1010110010;
    16'b0000000100100000: out_v[29] = 10'b0001000010;
    16'b1000000100000000: out_v[29] = 10'b1101100111;
    16'b0010000000000001: out_v[29] = 10'b1011100000;
    16'b0010000110000001: out_v[29] = 10'b1110100000;
    16'b0010110100000001: out_v[29] = 10'b0011110110;
    16'b1000000100000001: out_v[29] = 10'b1000100000;
    16'b1010000110000000: out_v[29] = 10'b1011111101;
    16'b0000000110100001: out_v[29] = 10'b0110011000;
    16'b1010010010100001: out_v[29] = 10'b1011110000;
    16'b0010000100000000: out_v[29] = 10'b1111100110;
    16'b1000010000100001: out_v[29] = 10'b0011000111;
    16'b1000010110100001: out_v[29] = 10'b0000100111;
    16'b0000010000100001: out_v[29] = 10'b1101000001;
    16'b0000000000100001: out_v[29] = 10'b0001001110;
    16'b0010000100100000: out_v[29] = 10'b1001110011;
    16'b1000010010100001: out_v[29] = 10'b0001000011;
    16'b1000000100100001: out_v[29] = 10'b1001001111;
    16'b1010010000100001: out_v[29] = 10'b1000111110;
    16'b0001010100100001: out_v[29] = 10'b1111001111;
    16'b0001010100000001: out_v[29] = 10'b0100010010;
    16'b0001010000000000: out_v[29] = 10'b0001001111;
    16'b0000010000000010: out_v[29] = 10'b0010110010;
    16'b0000010100000011: out_v[29] = 10'b1111110010;
    16'b0011010100100001: out_v[29] = 10'b0111100011;
    16'b0011010000100000: out_v[29] = 10'b0011100001;
    16'b1010000100100000: out_v[29] = 10'b1110011111;
    16'b1000000100100000: out_v[29] = 10'b1001000011;
    16'b1010000000000001: out_v[29] = 10'b0110100011;
    16'b1010000100100001: out_v[29] = 10'b1011101010;
    16'b1000000000100001: out_v[29] = 10'b1110100101;
    default: out_v[29] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000100100001: out_v[30] = 10'b0110000011;
    16'b0010000000000001: out_v[30] = 10'b0110001011;
    16'b0000000000100001: out_v[30] = 10'b0111011000;
    16'b0000010000000001: out_v[30] = 10'b1010101100;
    16'b0000000000000001: out_v[30] = 10'b1100111010;
    16'b0010010000000001: out_v[30] = 10'b1010111001;
    16'b0010000000000000: out_v[30] = 10'b0010100001;
    16'b0000010000100001: out_v[30] = 10'b1101000101;
    16'b0010000100000001: out_v[30] = 10'b1100011011;
    16'b0000000100000001: out_v[30] = 10'b1000111100;
    16'b0000001000000001: out_v[30] = 10'b1010101011;
    16'b0010010000000000: out_v[30] = 10'b1011000100;
    16'b0010001100000001: out_v[30] = 10'b0010101011;
    16'b0010001000000001: out_v[30] = 10'b0101010101;
    16'b0000001100000001: out_v[30] = 10'b1000101000;
    16'b0000010000000000: out_v[30] = 10'b1010100110;
    16'b0000000000000000: out_v[30] = 10'b0110101001;
    16'b0000010010100001: out_v[30] = 10'b1001011100;
    16'b0000001000000000: out_v[30] = 10'b0010111001;
    16'b0010010010100001: out_v[30] = 10'b1110111010;
    16'b0000000010100000: out_v[30] = 10'b0010110010;
    16'b0000000010000001: out_v[30] = 10'b0111110011;
    16'b0000000010000000: out_v[30] = 10'b1100010010;
    16'b0000010010100000: out_v[30] = 10'b0001011000;
    16'b0000000110000001: out_v[30] = 10'b0101101110;
    16'b0000000010100001: out_v[30] = 10'b0111000100;
    16'b0000010010000000: out_v[30] = 10'b0101010010;
    16'b0000000110000000: out_v[30] = 10'b0110110101;
    16'b0000010010000001: out_v[30] = 10'b1101011100;
    16'b0000010100000001: out_v[30] = 10'b0011010110;
    16'b0010000010100000: out_v[30] = 10'b1100100110;
    16'b0000000100000000: out_v[30] = 10'b1001110010;
    16'b0000010110000001: out_v[30] = 10'b0100000011;
    16'b0000001010100001: out_v[30] = 10'b1011000101;
    16'b0010010010100000: out_v[30] = 10'b0001111001;
    16'b0000001010100000: out_v[30] = 10'b0001010101;
    16'b0000011010100000: out_v[30] = 10'b0001011101;
    16'b0000011010100001: out_v[30] = 10'b1010111000;
    16'b0010011010100001: out_v[30] = 10'b0111100110;
    16'b0010000010100001: out_v[30] = 10'b0111110011;
    16'b0000011000000000: out_v[30] = 10'b1000100111;
    16'b0000011000000001: out_v[30] = 10'b0101010110;
    16'b0010010010000001: out_v[30] = 10'b0001111111;
    16'b0000011010000001: out_v[30] = 10'b0100000101;
    16'b0000011010100101: out_v[30] = 10'b0110010110;
    16'b0000000000100000: out_v[30] = 10'b0101010100;
    16'b0010011010100000: out_v[30] = 10'b0000110110;
    16'b0000010110100001: out_v[30] = 10'b1011000011;
    16'b0000000110100001: out_v[30] = 10'b0111101000;
    16'b0000011100000001: out_v[30] = 10'b1011001100;
    16'b0010010100000001: out_v[30] = 10'b1011110000;
    16'b0000010100000000: out_v[30] = 10'b0011011111;
    16'b0010010100000000: out_v[30] = 10'b1111111101;
    16'b0000010000100000: out_v[30] = 10'b0101010101;
    16'b0000010110100000: out_v[30] = 10'b1011001011;
    16'b0010010110100000: out_v[30] = 10'b1111100111;
    16'b0010010110100001: out_v[30] = 10'b1100011010;
    16'b0000010110000000: out_v[30] = 10'b0110000111;
    16'b0010000010000000: out_v[30] = 10'b1101001000;
    16'b0010010000000011: out_v[30] = 10'b1010001011;
    16'b0000010000000011: out_v[30] = 10'b1111110110;
    16'b0000010000000010: out_v[30] = 10'b1111000101;
    16'b0000010100010000: out_v[30] = 10'b1100100110;
    16'b0000000000010000: out_v[30] = 10'b1010011001;
    16'b0000010100010001: out_v[30] = 10'b1011011001;
    16'b0010010000000010: out_v[30] = 10'b1110011010;
    16'b0000010000010000: out_v[30] = 10'b1010000010;
    16'b0010000110100001: out_v[30] = 10'b0000101111;
    16'b0010010100100001: out_v[30] = 10'b0011000110;
    16'b0000010100100001: out_v[30] = 10'b1110100010;
    16'b0000001110100001: out_v[30] = 10'b1001100110;
    16'b0010010000100001: out_v[30] = 10'b0011000111;
    16'b0010000000100001: out_v[30] = 10'b1110110111;
    16'b0000011110100001: out_v[30] = 10'b0111111010;
    16'b0010010110000001: out_v[30] = 10'b0111001011;
    default: out_v[30] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010100001100000: out_v[31] = 10'b1001001101;
    16'b0000100000100000: out_v[31] = 10'b0000000111;
    16'b0010100000100000: out_v[31] = 10'b1000001111;
    16'b0010100000001000: out_v[31] = 10'b1000011101;
    16'b0000000000000000: out_v[31] = 10'b0010110011;
    16'b0010100000101000: out_v[31] = 10'b0101111100;
    16'b0000100001100000: out_v[31] = 10'b0110000011;
    16'b0010100000000000: out_v[31] = 10'b0101111110;
    16'b0010000000000000: out_v[31] = 10'b0101101000;
    16'b0000100000000000: out_v[31] = 10'b1111011101;
    16'b0000110010100000: out_v[31] = 10'b0010010101;
    16'b0000000000100000: out_v[31] = 10'b0010001101;
    16'b0000000001000000: out_v[31] = 10'b0111000101;
    16'b0000100000100010: out_v[31] = 10'b0111110011;
    16'b0000110000100000: out_v[31] = 10'b1001010110;
    16'b0010000001100000: out_v[31] = 10'b0001111011;
    16'b0000100000000010: out_v[31] = 10'b1000101011;
    16'b0000100000001000: out_v[31] = 10'b0001010100;
    16'b0000000001100000: out_v[31] = 10'b1001011011;
    16'b0010000000001000: out_v[31] = 10'b1011010010;
    16'b0010000000100000: out_v[31] = 10'b0001011011;
    16'b0000000000001000: out_v[31] = 10'b0011011101;
    16'b0010000000001010: out_v[31] = 10'b1010010110;
    16'b0000000001001000: out_v[31] = 10'b0010010101;
    16'b0000100001001000: out_v[31] = 10'b1100000011;
    16'b0010000000000010: out_v[31] = 10'b1001101010;
    16'b0000000000000010: out_v[31] = 10'b1001011000;
    16'b0100100000101000: out_v[31] = 10'b0111000001;
    16'b0010000000101000: out_v[31] = 10'b0110011100;
    16'b0100100000000000: out_v[31] = 10'b1111000000;
    16'b0000100000101000: out_v[31] = 10'b0111101100;
    16'b0110100000101000: out_v[31] = 10'b0001001011;
    16'b0000000000101000: out_v[31] = 10'b0110101000;
    16'b0010100000001010: out_v[31] = 10'b0110110101;
    16'b0110100000001000: out_v[31] = 10'b1101010100;
    16'b0010100000101010: out_v[31] = 10'b0110110010;
    16'b0010000001001000: out_v[31] = 10'b1000011100;
    16'b0100100000100000: out_v[31] = 10'b1111100110;
    16'b0000000001101000: out_v[31] = 10'b0000101010;
    16'b0010100001001000: out_v[31] = 10'b1010011010;
    16'b0000100101101000: out_v[31] = 10'b0010101110;
    16'b0000100001101000: out_v[31] = 10'b0011101001;
    16'b0010100001101000: out_v[31] = 10'b0110011011;
    16'b0010000001101000: out_v[31] = 10'b1111001011;
    16'b0010000001000000: out_v[31] = 10'b1110101000;
    16'b0000100101001000: out_v[31] = 10'b1001100110;
    16'b0000000101001000: out_v[31] = 10'b0111010000;
    16'b0010000100001000: out_v[31] = 10'b1011100000;
    16'b0010100101001000: out_v[31] = 10'b0101001110;
    16'b0010100100001000: out_v[31] = 10'b1110100110;
    16'b0010110010101000: out_v[31] = 10'b0011010011;
    16'b0010000101001000: out_v[31] = 10'b0001011111;
    16'b0000000000001001: out_v[31] = 10'b1110111000;
    16'b0000100000001001: out_v[31] = 10'b0100100010;
    16'b0000100001000000: out_v[31] = 10'b0110100000;
    16'b0000000000001010: out_v[31] = 10'b1011101000;
    16'b0000100000000001: out_v[31] = 10'b0000111000;
    16'b0000100000001010: out_v[31] = 10'b0000111111;
    16'b0000100000101010: out_v[31] = 10'b0001000010;
    16'b0000100101000000: out_v[31] = 10'b0001111100;
    16'b0000100000101001: out_v[31] = 10'b1011100111;
    16'b0000000000000001: out_v[31] = 10'b0001111111;
    16'b0010100000100010: out_v[31] = 10'b0100110011;
    16'b0001100000101000: out_v[31] = 10'b0001000010;
    16'b0011100000100000: out_v[31] = 10'b0011011001;
    16'b0011100000101000: out_v[31] = 10'b1111101011;
    16'b0110100000100000: out_v[31] = 10'b0010111111;
    16'b0001100000001000: out_v[31] = 10'b1010100100;
    16'b0011100000001000: out_v[31] = 10'b1101100111;
    16'b0010000010001000: out_v[31] = 10'b1111001011;
    16'b0010100100000000: out_v[31] = 10'b1110010100;
    16'b0010100101101000: out_v[31] = 10'b1010001000;
    16'b0010100111001000: out_v[31] = 10'b1001111111;
    16'b0010110111001000: out_v[31] = 10'b0010011111;
    16'b0000000100001000: out_v[31] = 10'b1111000001;
    16'b0010100101100000: out_v[31] = 10'b1110110110;
    16'b0010100010001000: out_v[31] = 10'b1010000101;
    16'b0010100101000000: out_v[31] = 10'b1111010011;
    16'b0010100000001001: out_v[31] = 10'b1000010101;
    16'b0010100001000000: out_v[31] = 10'b1001110111;
    16'b0010000000001001: out_v[31] = 10'b0111111010;
    16'b0010000000000001: out_v[31] = 10'b1100101011;
    16'b0010010010101000: out_v[31] = 10'b1001001011;
    default: out_v[31] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1101100000000010: out_v[32] = 10'b1010011111;
    16'b1101101011000010: out_v[32] = 10'b1001001001;
    16'b0100101011000000: out_v[32] = 10'b1010100111;
    16'b1001100000000000: out_v[32] = 10'b0100100011;
    16'b1001101011000010: out_v[32] = 10'b1010011111;
    16'b1101100001000010: out_v[32] = 10'b1101111110;
    16'b1000101011000000: out_v[32] = 10'b0111000111;
    16'b1001101000000010: out_v[32] = 10'b1101010100;
    16'b1101100000010010: out_v[32] = 10'b1110111010;
    16'b1101100010000010: out_v[32] = 10'b0111100110;
    16'b1101101011000000: out_v[32] = 10'b0111101111;
    16'b1100101011000010: out_v[32] = 10'b0011010101;
    16'b1100101011000000: out_v[32] = 10'b0101100110;
    16'b0001100000000000: out_v[32] = 10'b0010011011;
    16'b1101100011000000: out_v[32] = 10'b0010011101;
    16'b1101100011000010: out_v[32] = 10'b1101000110;
    16'b1000101010000010: out_v[32] = 10'b0100000111;
    16'b1000101011000010: out_v[32] = 10'b1010110011;
    16'b1001100000000010: out_v[32] = 10'b1100001001;
    16'b0101100000010010: out_v[32] = 10'b1011111110;
    16'b0100101011000010: out_v[32] = 10'b0111110110;
    16'b0001100000010010: out_v[32] = 10'b0001110111;
    16'b1101100011010010: out_v[32] = 10'b1111011110;
    16'b1000101010000000: out_v[32] = 10'b1110000111;
    16'b1001100001000000: out_v[32] = 10'b1100001011;
    16'b1101100001000000: out_v[32] = 10'b1110110001;
    16'b1101101011010010: out_v[32] = 10'b1001001110;
    16'b1001000000000010: out_v[32] = 10'b0010110011;
    16'b0100101011010000: out_v[32] = 10'b1111110101;
    16'b1101100000000000: out_v[32] = 10'b1011110011;
    16'b1100101010000000: out_v[32] = 10'b1010111011;
    16'b1101100001010010: out_v[32] = 10'b0111101010;
    16'b1101101010000000: out_v[32] = 10'b1110110111;
    16'b1100101010000010: out_v[32] = 10'b0001010011;
    16'b1001100000010010: out_v[32] = 10'b1001101110;
    16'b0100101011010010: out_v[32] = 10'b1011000011;
    16'b1101101010000010: out_v[32] = 10'b1011001101;
    16'b1100001011000010: out_v[32] = 10'b1110011001;
    16'b1001110000000010: out_v[32] = 10'b0110101001;
    16'b1100001011000000: out_v[32] = 10'b1011110011;
    16'b0000110000000010: out_v[32] = 10'b1011100110;
    16'b0001010000000010: out_v[32] = 10'b1100001001;
    16'b0000000000000000: out_v[32] = 10'b1011100111;
    16'b0001000000000000: out_v[32] = 10'b1111100110;
    16'b0001001000000010: out_v[32] = 10'b0100001111;
    16'b0000000000000010: out_v[32] = 10'b1001101011;
    16'b0001001000000000: out_v[32] = 10'b1001011011;
    16'b0001011000000000: out_v[32] = 10'b0010010111;
    16'b0000100000000010: out_v[32] = 10'b1000101111;
    16'b1000110000000010: out_v[32] = 10'b0011001010;
    16'b0001011000000010: out_v[32] = 10'b0011010010;
    16'b0000010000000010: out_v[32] = 10'b1011110001;
    16'b0001000000000010: out_v[32] = 10'b0111001000;
    16'b0001110000000010: out_v[32] = 10'b1111100010;
    16'b1000100000000010: out_v[32] = 10'b1111101000;
    16'b1000110000000000: out_v[32] = 10'b1100100110;
    16'b0001010000000000: out_v[32] = 10'b1001111001;
    16'b1001110000000000: out_v[32] = 10'b1111000100;
    16'b0001010010000010: out_v[32] = 10'b0010010011;
    16'b0000011010000010: out_v[32] = 10'b0101001101;
    16'b1001111010000010: out_v[32] = 10'b1010011000;
    16'b1001110010000010: out_v[32] = 10'b0100010111;
    16'b1001010000000010: out_v[32] = 10'b0111100110;
    16'b1101010000000010: out_v[32] = 10'b1101000111;
    16'b1001110010000000: out_v[32] = 10'b1001000100;
    16'b0000001010000010: out_v[32] = 10'b1100011101;
    16'b1001110011000010: out_v[32] = 10'b0011011100;
    16'b1001010010000010: out_v[32] = 10'b0000110010;
    16'b1001110010010010: out_v[32] = 10'b1111011011;
    16'b1001100010010000: out_v[32] = 10'b0011011000;
    16'b1001100010000000: out_v[32] = 10'b1011100110;
    16'b1100010000000010: out_v[32] = 10'b1001101111;
    16'b1000111010000010: out_v[32] = 10'b1101001000;
    16'b1001111000000000: out_v[32] = 10'b1001101100;
    16'b1101110000000010: out_v[32] = 10'b0011100111;
    16'b1001110011000000: out_v[32] = 10'b0010111110;
    16'b1101010010000010: out_v[32] = 10'b0111010110;
    16'b1001111010000000: out_v[32] = 10'b1011011011;
    16'b0001000010000010: out_v[32] = 10'b0010111111;
    16'b0001011010000010: out_v[32] = 10'b1000100111;
    16'b1101110000000000: out_v[32] = 10'b1100110101;
    16'b1001100010000010: out_v[32] = 10'b1011110110;
    16'b1001110010010000: out_v[32] = 10'b1001100011;
    16'b1000110010000000: out_v[32] = 10'b1110000100;
    16'b1101110010000000: out_v[32] = 10'b1010110010;
    16'b1001000010000010: out_v[32] = 10'b1111000000;
    16'b1101000000000010: out_v[32] = 10'b1110010010;
    16'b0001110010000000: out_v[32] = 10'b0001011111;
    16'b1000111010000000: out_v[32] = 10'b0011001010;
    16'b1101110010000010: out_v[32] = 10'b0111110011;
    16'b1000010000000010: out_v[32] = 10'b1000100101;
    16'b0001111000000010: out_v[32] = 10'b0110001101;
    16'b1000011010000010: out_v[32] = 10'b1010011011;
    16'b0101011010000010: out_v[32] = 10'b1111011011;
    16'b0000011000000010: out_v[32] = 10'b0100011101;
    16'b0100011010000010: out_v[32] = 10'b0100001010;
    16'b0110011010000010: out_v[32] = 10'b1010100011;
    16'b0001110000000000: out_v[32] = 10'b1101011001;
    16'b0001110000010000: out_v[32] = 10'b1011011001;
    16'b1001110000010000: out_v[32] = 10'b0110001011;
    16'b0000111010000010: out_v[32] = 10'b0110111010;
    16'b0010011010000010: out_v[32] = 10'b0001111010;
    16'b0110111010000010: out_v[32] = 10'b0011011100;
    16'b0101111010000010: out_v[32] = 10'b1100001010;
    16'b1001110000010010: out_v[32] = 10'b1010001001;
    16'b0000101010000010: out_v[32] = 10'b1001001101;
    16'b1100111010000010: out_v[32] = 10'b1100101111;
    16'b0001100000000010: out_v[32] = 10'b0111101000;
    16'b1100011010000010: out_v[32] = 10'b1011101011;
    16'b0001110000010010: out_v[32] = 10'b1010100100;
    16'b1101111010000010: out_v[32] = 10'b1110001110;
    16'b0100111010000010: out_v[32] = 10'b0011000111;
    16'b0001111010000010: out_v[32] = 10'b0011111010;
    16'b0100001010000010: out_v[32] = 10'b0011011100;
    16'b0000011010000000: out_v[32] = 10'b0111100101;
    16'b0000001000000010: out_v[32] = 10'b1101001101;
    16'b0100111010000000: out_v[32] = 10'b1001101011;
    16'b0000111010000000: out_v[32] = 10'b1100011000;
    16'b0001111000000000: out_v[32] = 10'b1100001001;
    16'b0000111000000000: out_v[32] = 10'b1000011010;
    16'b1100001010000010: out_v[32] = 10'b1111011110;
    16'b0100111010010010: out_v[32] = 10'b1001001010;
    16'b0100011010000000: out_v[32] = 10'b0110101000;
    16'b0001111001000000: out_v[32] = 10'b0010011011;
    16'b0001011001000010: out_v[32] = 10'b0100011101;
    16'b0000010000000000: out_v[32] = 10'b1010101100;
    16'b0001110001000010: out_v[32] = 10'b1101001101;
    16'b0000110000000000: out_v[32] = 10'b1010010000;
    16'b0001110001000000: out_v[32] = 10'b1000011010;
    16'b0001010001000000: out_v[32] = 10'b0100011011;
    16'b0001011001000000: out_v[32] = 10'b1111001011;
    16'b0001101001000000: out_v[32] = 10'b0101011110;
    16'b0001111001000010: out_v[32] = 10'b1011010100;
    16'b0000111001000000: out_v[32] = 10'b0011101111;
    16'b0000010011000010: out_v[32] = 10'b1101010010;
    16'b0000110001000000: out_v[32] = 10'b1000010010;
    16'b0000110011000000: out_v[32] = 10'b0110001011;
    16'b0000110010000000: out_v[32] = 10'b0100011010;
    16'b0001010001000010: out_v[32] = 10'b1001111001;
    16'b0000010010000010: out_v[32] = 10'b1100010101;
    16'b0101110001000000: out_v[32] = 10'b1000111010;
    16'b0100011011000000: out_v[32] = 10'b0010110101;
    16'b0100111011000000: out_v[32] = 10'b0111010010;
    16'b0000111011000010: out_v[32] = 10'b0101100110;
    16'b0001101001000010: out_v[32] = 10'b0001100100;
    16'b0100001011000000: out_v[32] = 10'b0011100111;
    16'b1001010000000000: out_v[32] = 10'b0111001000;
    16'b0000001000000000: out_v[32] = 10'b0010100111;
    16'b0000011011000000: out_v[32] = 10'b0011100111;
    16'b0001101000000010: out_v[32] = 10'b1101100000;
    16'b0100111011000010: out_v[32] = 10'b1001100110;
    16'b1001000000000000: out_v[32] = 10'b1011000110;
    16'b0100001010000000: out_v[32] = 10'b1000110011;
    16'b0000001011000000: out_v[32] = 10'b0010110110;
    16'b1100011011000000: out_v[32] = 10'b0010011110;
    16'b0001100001000010: out_v[32] = 10'b1011110010;
    16'b1000011011000000: out_v[32] = 10'b1001111011;
    16'b0000011000000000: out_v[32] = 10'b1001100101;
    16'b0000001010000000: out_v[32] = 10'b1001001010;
    16'b1100011010000000: out_v[32] = 10'b1110100110;
    16'b0000111011000000: out_v[32] = 10'b0011001110;
    16'b0101011010000000: out_v[32] = 10'b1001111011;
    16'b1101010010000000: out_v[32] = 10'b0010100111;
    16'b0101010011000000: out_v[32] = 10'b1100001001;
    16'b0001010011100000: out_v[32] = 10'b1111101011;
    16'b1101011011000000: out_v[32] = 10'b0001010011;
    16'b1001010011000000: out_v[32] = 10'b1111010010;
    16'b0101010010100000: out_v[32] = 10'b1110101111;
    16'b1101010011100000: out_v[32] = 10'b1100001011;
    16'b1101010011000000: out_v[32] = 10'b0111101100;
    16'b0101011011000000: out_v[32] = 10'b1010100001;
    16'b0101010011100000: out_v[32] = 10'b1010110011;
    16'b0101000010000000: out_v[32] = 10'b1110110111;
    16'b1001010011100000: out_v[32] = 10'b0111111111;
    16'b0101010000000000: out_v[32] = 10'b1001101101;
    16'b0101010010000000: out_v[32] = 10'b1110101101;
    16'b1101010000000000: out_v[32] = 10'b1011111011;
    16'b1101010001000000: out_v[32] = 10'b0111110010;
    16'b1101000000000000: out_v[32] = 10'b1011010010;
    16'b0001011010000000: out_v[32] = 10'b0101000001;
    16'b0001010010100000: out_v[32] = 10'b1111101011;
    16'b1001010000000011: out_v[32] = 10'b1011011010;
    16'b1101010010100000: out_v[32] = 10'b0111101001;
    16'b1101011010000000: out_v[32] = 10'b1010110111;
    16'b1101000010000000: out_v[32] = 10'b1010011100;
    16'b0001010000100000: out_v[32] = 10'b1111101001;
    16'b0101010000100000: out_v[32] = 10'b1111111110;
    16'b1101010001100000: out_v[32] = 10'b1000111111;
    16'b0001010011000000: out_v[32] = 10'b1111011011;
    16'b0001010010000000: out_v[32] = 10'b1111010011;
    16'b1001010010000000: out_v[32] = 10'b1110110001;
    16'b1101010000000011: out_v[32] = 10'b1111000110;
    16'b0011011001000010: out_v[32] = 10'b0101100111;
    16'b0011011000000010: out_v[32] = 10'b0111110010;
    16'b0011111000000010: out_v[32] = 10'b1010101011;
    16'b0001000001000010: out_v[32] = 10'b1001101011;
    16'b0011111001000010: out_v[32] = 10'b0101111011;
    16'b0011110000000010: out_v[32] = 10'b1111001001;
    16'b0000110001000010: out_v[32] = 10'b1010001101;
    16'b0011110001000010: out_v[32] = 10'b1101110101;
    16'b0011100001000010: out_v[32] = 10'b0100111111;
    16'b0001001001000010: out_v[32] = 10'b1010101101;
    16'b0011100000000010: out_v[32] = 10'b1100100001;
    16'b0011010000000010: out_v[32] = 10'b1111100101;
    16'b0011101001000010: out_v[32] = 10'b1101011010;
    16'b1000111000000000: out_v[32] = 10'b0101011110;
    16'b1001110001000010: out_v[32] = 10'b0111110010;
    16'b1000010000000000: out_v[32] = 10'b0000100111;
    16'b0001111011000000: out_v[32] = 10'b1111000010;
    16'b1001110001000000: out_v[32] = 10'b0111110010;
    16'b1100111011000010: out_v[32] = 10'b0100110010;
    16'b1001111000000010: out_v[32] = 10'b1000101111;
    16'b1001111001000000: out_v[32] = 10'b1000010011;
    16'b0001101000000000: out_v[32] = 10'b0000110101;
    16'b1000111011000000: out_v[32] = 10'b0111010001;
    16'b0001111011000010: out_v[32] = 10'b1100010011;
    16'b1100111011000000: out_v[32] = 10'b0110111011;
    16'b1001111001000010: out_v[32] = 10'b1011101010;
    16'b1001011000000000: out_v[32] = 10'b1101100010;
    16'b1000111011000010: out_v[32] = 10'b0101110111;
    16'b0000011011000010: out_v[32] = 10'b1111000001;
    16'b0000011001000010: out_v[32] = 10'b0101001100;
    16'b0000111001000010: out_v[32] = 10'b0001110101;
    default: out_v[32] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010000010010000: out_v[33] = 10'b0010110011;
    16'b0010100010000000: out_v[33] = 10'b0111000001;
    16'b0011100010000000: out_v[33] = 10'b0101100011;
    16'b0010000010000000: out_v[33] = 10'b0011011101;
    16'b0011000010000000: out_v[33] = 10'b0010110101;
    16'b0011100000000000: out_v[33] = 10'b1011001011;
    16'b0001000000010000: out_v[33] = 10'b0110010111;
    16'b0010000000000000: out_v[33] = 10'b0011001101;
    16'b0000000010010000: out_v[33] = 10'b1101100011;
    16'b0010100010010000: out_v[33] = 10'b0101100011;
    16'b0000100010010000: out_v[33] = 10'b1001100111;
    16'b0010000000010000: out_v[33] = 10'b1000011000;
    16'b0000000000010000: out_v[33] = 10'b1101100111;
    16'b0000100000000000: out_v[33] = 10'b0011011011;
    16'b0000000010000000: out_v[33] = 10'b1000000100;
    16'b0000100000010000: out_v[33] = 10'b0101000101;
    16'b0000100010000000: out_v[33] = 10'b0010110010;
    16'b0010100000000000: out_v[33] = 10'b1010001000;
    16'b0001000010010000: out_v[33] = 10'b0010011111;
    16'b0011100010010000: out_v[33] = 10'b0111111010;
    16'b0001000010000000: out_v[33] = 10'b0111001001;
    16'b0000000000000000: out_v[33] = 10'b1010011001;
    16'b0010100000010000: out_v[33] = 10'b1100001100;
    16'b0010100000010010: out_v[33] = 10'b0010111001;
    16'b0010100000000110: out_v[33] = 10'b1011010000;
    16'b0010100000010110: out_v[33] = 10'b0011011010;
    16'b0000100000010110: out_v[33] = 10'b1001100111;
    16'b0010100000000010: out_v[33] = 10'b0011100111;
    16'b0000100000010010: out_v[33] = 10'b0001010110;
    16'b0000000000010110: out_v[33] = 10'b0101110001;
    16'b0010000000010110: out_v[33] = 10'b1001010100;
    16'b0010000000010010: out_v[33] = 10'b1000011111;
    16'b0000000000010100: out_v[33] = 10'b1101111010;
    16'b0010000000000010: out_v[33] = 10'b1011100110;
    16'b0010101000000000: out_v[33] = 10'b0000001101;
    16'b0000100010010110: out_v[33] = 10'b1000101011;
    16'b0000000000010010: out_v[33] = 10'b1010100101;
    16'b0000000010010110: out_v[33] = 10'b0000001010;
    16'b0010000000010100: out_v[33] = 10'b1011110011;
    16'b0001100010000000: out_v[33] = 10'b1100100100;
    16'b0001100000000000: out_v[33] = 10'b1100100010;
    16'b0001000000000000: out_v[33] = 10'b0001110000;
    16'b0000100000000100: out_v[33] = 10'b1010110001;
    16'b1010000000010000: out_v[33] = 10'b1001100111;
    default: out_v[33] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001000000000000: out_v[34] = 10'b0111111101;
    16'b0001000000110000: out_v[34] = 10'b1000110011;
    16'b0000000000110000: out_v[34] = 10'b1000000011;
    16'b0001000000010000: out_v[34] = 10'b0000010000;
    16'b0001000000100000: out_v[34] = 10'b1010011000;
    16'b0000000000100000: out_v[34] = 10'b0010011011;
    16'b0000000000010000: out_v[34] = 10'b0110110001;
    16'b0000000001010100: out_v[34] = 10'b0110110010;
    16'b0000000000010100: out_v[34] = 10'b0011110011;
    16'b0000000000000000: out_v[34] = 10'b1101110011;
    16'b0000000001110000: out_v[34] = 10'b1100011101;
    16'b0001000001110100: out_v[34] = 10'b0001011111;
    16'b0001000001100000: out_v[34] = 10'b0101011010;
    16'b0001000001010000: out_v[34] = 10'b0011011111;
    16'b0000000001110100: out_v[34] = 10'b0100001111;
    16'b0000000001100100: out_v[34] = 10'b1010001100;
    16'b0001000000110100: out_v[34] = 10'b0100111101;
    16'b0001000010110000: out_v[34] = 10'b1011010011;
    16'b0000000000110100: out_v[34] = 10'b0101000011;
    16'b0000000000100100: out_v[34] = 10'b0000011101;
    16'b0000000001000100: out_v[34] = 10'b1000111100;
    16'b0001000010100000: out_v[34] = 10'b0010110001;
    16'b0000000000000100: out_v[34] = 10'b1110100101;
    16'b0001000001110000: out_v[34] = 10'b1110011111;
    16'b0001000010010000: out_v[34] = 10'b0101010100;
    16'b0000000001010000: out_v[34] = 10'b0011001010;
    16'b0000000010100000: out_v[34] = 10'b1100101100;
    16'b0000000001000000: out_v[34] = 10'b1001000011;
    16'b0000000010000000: out_v[34] = 10'b0110010000;
    16'b0000000001000101: out_v[34] = 10'b0011110010;
    16'b0001000001000100: out_v[34] = 10'b1100000000;
    16'b0001000001000000: out_v[34] = 10'b1011001011;
    16'b0000000001100101: out_v[34] = 10'b0100100110;
    16'b0001000000100100: out_v[34] = 10'b1111110100;
    16'b0001000001100100: out_v[34] = 10'b1101000110;
    16'b0001000000100101: out_v[34] = 10'b0011000110;
    16'b0000000001100000: out_v[34] = 10'b1100110101;
    16'b0001000010000000: out_v[34] = 10'b1100011111;
    16'b0001000001100101: out_v[34] = 10'b0010110100;
    16'b0001000000000100: out_v[34] = 10'b1110100101;
    16'b0000000000100101: out_v[34] = 10'b1000100111;
    16'b0000000000100001: out_v[34] = 10'b1011010011;
    16'b0001000000100001: out_v[34] = 10'b0100111110;
    16'b0000000000000101: out_v[34] = 10'b0010101111;
    16'b0001000000000101: out_v[34] = 10'b1010011110;
    16'b0000000000000001: out_v[34] = 10'b1010110100;
    16'b0001000000000001: out_v[34] = 10'b1101000110;
    16'b0010000000100000: out_v[34] = 10'b0001101010;
    16'b0001000001010100: out_v[34] = 10'b0001000101;
    16'b0001000000010100: out_v[34] = 10'b1001001000;
    16'b0011000000100000: out_v[34] = 10'b0111001001;
    16'b0001010000010000: out_v[34] = 10'b1111001010;
    16'b0001010000110000: out_v[34] = 10'b0111110100;
    16'b0001001000010000: out_v[34] = 10'b1110110000;
    16'b0000100000100000: out_v[34] = 10'b0111001111;
    16'b0000100000110000: out_v[34] = 10'b1011011111;
    16'b0001001010000000: out_v[34] = 10'b1100110001;
    16'b0000001000100000: out_v[34] = 10'b1001100000;
    16'b0001010000000000: out_v[34] = 10'b0111110110;
    16'b0001010000100000: out_v[34] = 10'b0011000010;
    16'b0000010000100000: out_v[34] = 10'b0001101111;
    16'b0010000000000000: out_v[34] = 10'b1001101001;
    16'b0011000000110000: out_v[34] = 10'b1011001110;
    16'b0010000000110000: out_v[34] = 10'b1011001011;
    16'b0011000000000000: out_v[34] = 10'b1100010111;
    16'b0000010000000000: out_v[34] = 10'b1110101000;
    16'b0000010000010000: out_v[34] = 10'b1101100011;
    16'b0011000000010000: out_v[34] = 10'b1010011101;
    16'b0010000000010000: out_v[34] = 10'b0101100101;
    16'b0000010000110000: out_v[34] = 10'b0010100110;
    default: out_v[34] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000000000000: out_v[35] = 10'b0101110110;
    16'b0000000100000000: out_v[35] = 10'b0100110011;
    16'b1000001100000000: out_v[35] = 10'b0010110010;
    16'b0000001000000000: out_v[35] = 10'b1110001001;
    16'b1000000000000000: out_v[35] = 10'b0010011100;
    16'b1000001000000000: out_v[35] = 10'b1101110100;
    16'b0000001001000000: out_v[35] = 10'b1110010000;
    16'b0000000000000001: out_v[35] = 10'b0000001100;
    16'b0000001100000000: out_v[35] = 10'b0110001000;
    16'b0000000100000001: out_v[35] = 10'b1000001010;
    16'b1000001000000010: out_v[35] = 10'b1111100011;
    16'b0000000110000001: out_v[35] = 10'b0111010001;
    16'b1000001001000000: out_v[35] = 10'b0110110001;
    16'b0000001000000010: out_v[35] = 10'b1100000111;
    16'b0000001000000001: out_v[35] = 10'b0001000101;
    16'b0000000010000001: out_v[35] = 10'b0100100101;
    16'b0000000010000000: out_v[35] = 10'b0001001011;
    16'b1000000000000010: out_v[35] = 10'b0010001100;
    16'b0000000000000010: out_v[35] = 10'b0000000101;
    16'b1000000000000001: out_v[35] = 10'b0000001110;
    16'b1000000100000000: out_v[35] = 10'b1100001010;
    16'b1000000010000001: out_v[35] = 10'b1010101000;
    16'b1000000110000001: out_v[35] = 10'b1001011111;
    16'b0000000110000000: out_v[35] = 10'b0110100001;
    16'b1000000100000001: out_v[35] = 10'b1011111111;
    16'b1000000110000000: out_v[35] = 10'b0000011001;
    16'b0000000001000000: out_v[35] = 10'b0011001010;
    16'b0000000000100000: out_v[35] = 10'b1111000000;
    16'b0000001101000000: out_v[35] = 10'b0011101001;
    default: out_v[35] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1000000000000000: out_v[36] = 10'b1000110111;
    16'b0101000000000100: out_v[36] = 10'b1001010111;
    16'b1001000000000100: out_v[36] = 10'b0011100111;
    16'b0000000000000000: out_v[36] = 10'b0010101101;
    16'b0000001000000000: out_v[36] = 10'b1101100100;
    16'b0100001000000000: out_v[36] = 10'b1010001001;
    16'b0100000000000000: out_v[36] = 10'b0011011011;
    16'b0101000000000000: out_v[36] = 10'b1010001001;
    16'b0000000000000100: out_v[36] = 10'b1011011110;
    16'b1100000000100000: out_v[36] = 10'b0001000011;
    16'b0100001000100000: out_v[36] = 10'b1000110101;
    16'b1100000000000100: out_v[36] = 10'b1011011011;
    16'b1100000000000000: out_v[36] = 10'b1100100011;
    16'b0001000000000000: out_v[36] = 10'b1101110011;
    16'b0001000000000100: out_v[36] = 10'b0100110011;
    16'b0100000000100000: out_v[36] = 10'b0100101111;
    16'b1000001000000000: out_v[36] = 10'b1100110011;
    16'b1001000000000000: out_v[36] = 10'b1001110111;
    16'b0101010000000100: out_v[36] = 10'b0011101011;
    16'b1100001000000000: out_v[36] = 10'b0101010101;
    16'b0000000000100000: out_v[36] = 10'b0101001010;
    16'b0001010000000100: out_v[36] = 10'b0000110011;
    16'b0100000000000100: out_v[36] = 10'b0000011101;
    16'b1101000000000100: out_v[36] = 10'b0111011010;
    16'b1101010000000100: out_v[36] = 10'b0011111111;
    16'b1100001000100000: out_v[36] = 10'b0001110001;
    16'b0000010000000100: out_v[36] = 10'b1110100101;
    16'b1000000000000100: out_v[36] = 10'b0001100110;
    16'b0100010000000100: out_v[36] = 10'b1001001111;
    16'b0000001000100000: out_v[36] = 10'b0001010110;
    16'b1101000000000000: out_v[36] = 10'b0001110110;
    16'b1001010000000100: out_v[36] = 10'b0110011001;
    16'b0100010000000000: out_v[36] = 10'b0011110011;
    16'b0000010000000000: out_v[36] = 10'b1100000111;
    16'b0100001000000100: out_v[36] = 10'b0010011100;
    16'b0000001000100100: out_v[36] = 10'b1001000011;
    16'b1100000000100100: out_v[36] = 10'b0100011100;
    16'b0000001000000100: out_v[36] = 10'b0100101100;
    16'b0100000000100100: out_v[36] = 10'b1100110110;
    16'b0101001000100100: out_v[36] = 10'b0100011000;
    16'b1000001000000100: out_v[36] = 10'b0111100100;
    16'b1000001000100100: out_v[36] = 10'b0000011010;
    16'b0101000000100100: out_v[36] = 10'b1101000001;
    16'b0101001000000100: out_v[36] = 10'b1001011001;
    16'b0101001000000000: out_v[36] = 10'b1100100000;
    16'b0001001000000100: out_v[36] = 10'b1111011010;
    16'b1000000000100100: out_v[36] = 10'b0010110101;
    16'b0100001000100100: out_v[36] = 10'b1100000110;
    16'b1000001000100000: out_v[36] = 10'b1111001101;
    16'b0000000000100100: out_v[36] = 10'b0111110100;
    16'b0001001000000000: out_v[36] = 10'b0011000101;
    16'b1000000000100000: out_v[36] = 10'b1111001100;
    16'b0001001000100000: out_v[36] = 10'b1001110101;
    16'b1001001000000100: out_v[36] = 10'b0111010110;
    16'b0000011000000100: out_v[36] = 10'b0011001111;
    16'b0100011000000000: out_v[36] = 10'b1011000000;
    16'b0100011000100000: out_v[36] = 10'b0011010011;
    16'b0100010000100000: out_v[36] = 10'b0111110001;
    16'b0100011000000100: out_v[36] = 10'b0001110111;
    16'b0101011000000100: out_v[36] = 10'b1100100001;
    16'b0100010000100100: out_v[36] = 10'b1001001011;
    16'b0100011000100100: out_v[36] = 10'b0111001101;
    16'b0101011000100100: out_v[36] = 10'b0100110010;
    16'b0000011000100100: out_v[36] = 10'b0101001110;
    16'b0000011000100000: out_v[36] = 10'b0000010000;
    16'b0101001000100000: out_v[36] = 10'b0011110010;
    16'b0101011000100000: out_v[36] = 10'b1101000101;
    16'b0001001000100100: out_v[36] = 10'b0110011010;
    16'b0001011000000000: out_v[36] = 10'b1100010011;
    16'b0001011000100000: out_v[36] = 10'b0100100010;
    16'b0101011000000000: out_v[36] = 10'b0111111001;
    16'b1000011000100000: out_v[36] = 10'b1011100101;
    16'b1001011000100000: out_v[36] = 10'b0111111001;
    16'b1000011000000000: out_v[36] = 10'b0110011010;
    16'b1001001000100000: out_v[36] = 10'b1100110000;
    16'b1001001000000000: out_v[36] = 10'b0000110111;
    16'b0000011000000000: out_v[36] = 10'b1000101000;
    16'b1000011000100100: out_v[36] = 10'b1010111111;
    16'b1000010000000100: out_v[36] = 10'b0110111001;
    16'b0000010000100000: out_v[36] = 10'b0111100011;
    16'b1001011000000100: out_v[36] = 10'b1101001010;
    16'b0001000000100100: out_v[36] = 10'b1111100010;
    16'b0101010000000000: out_v[36] = 10'b0011100111;
    16'b0001010000000000: out_v[36] = 10'b0010101010;
    16'b0001011000100100: out_v[36] = 10'b1000101110;
    16'b0001010000100000: out_v[36] = 10'b1111001010;
    16'b1000010000100000: out_v[36] = 10'b1001010011;
    16'b0101010000100000: out_v[36] = 10'b0110100010;
    16'b0001011000000100: out_v[36] = 10'b1110100001;
    16'b0001010000100100: out_v[36] = 10'b0110110011;
    default: out_v[36] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001000000000110: out_v[37] = 10'b0011111000;
    16'b1001010010000010: out_v[37] = 10'b0011011011;
    16'b1001010010110110: out_v[37] = 10'b1011001110;
    16'b1001010010010110: out_v[37] = 10'b0101110110;
    16'b0001000010000110: out_v[37] = 10'b1010100101;
    16'b1001000000000010: out_v[37] = 10'b1101000000;
    16'b1001000010110010: out_v[37] = 10'b1001011111;
    16'b1000010010010110: out_v[37] = 10'b1101100001;
    16'b1001010010110010: out_v[37] = 10'b1011010001;
    16'b1001010010010010: out_v[37] = 10'b0011110111;
    16'b1001000000100010: out_v[37] = 10'b1100100111;
    16'b1001010010000110: out_v[37] = 10'b0000100100;
    16'b0001010010000110: out_v[37] = 10'b1011100010;
    16'b0000010010000110: out_v[37] = 10'b0001001001;
    16'b1000010010110010: out_v[37] = 10'b1011010011;
    16'b1001000000000110: out_v[37] = 10'b0010110111;
    16'b1001000010000110: out_v[37] = 10'b0011100110;
    16'b1001000010000100: out_v[37] = 10'b1000111111;
    16'b1000010010110110: out_v[37] = 10'b0100110011;
    16'b1001000010000010: out_v[37] = 10'b0011010000;
    16'b0000010010010110: out_v[37] = 10'b1001111010;
    16'b1001010010100010: out_v[37] = 10'b0111000100;
    16'b1000010010010100: out_v[37] = 10'b1000100101;
    16'b1001000000110010: out_v[37] = 10'b1101100110;
    16'b1001000000100000: out_v[37] = 10'b0011011011;
    16'b0001000000000100: out_v[37] = 10'b1101001011;
    16'b0001000010000100: out_v[37] = 10'b0010101011;
    16'b0001010010000100: out_v[37] = 10'b0001111001;
    16'b1011010010110110: out_v[37] = 10'b1111111111;
    16'b1001000010100010: out_v[37] = 10'b1101010110;
    16'b1011010010010110: out_v[37] = 10'b0110110100;
    16'b1000010010010010: out_v[37] = 10'b0101100001;
    16'b1001010010110000: out_v[37] = 10'b0111010111;
    16'b0001010010100110: out_v[37] = 10'b1100101001;
    16'b0001010010010110: out_v[37] = 10'b1110000010;
    16'b1001000010100110: out_v[37] = 10'b1000111011;
    16'b0000010010010100: out_v[37] = 10'b0010011011;
    16'b1001000010010110: out_v[37] = 10'b0011011101;
    16'b1001000010010010: out_v[37] = 10'b1011010111;
    16'b1001000000000100: out_v[37] = 10'b1100011110;
    16'b1000010010000110: out_v[37] = 10'b1111100110;
    16'b1001010010000100: out_v[37] = 10'b1000110001;
    16'b1001010010100110: out_v[37] = 10'b0010011011;
    16'b1001000000100110: out_v[37] = 10'b1001101011;
    16'b0000010010000100: out_v[37] = 10'b1101110010;
    16'b0001010010000010: out_v[37] = 10'b0100111111;
    16'b0000010010110110: out_v[37] = 10'b1011010111;
    16'b0001000010000010: out_v[37] = 10'b0000110001;
    16'b0010010000010110: out_v[37] = 10'b1111111110;
    16'b0000000000100000: out_v[37] = 10'b0001100011;
    16'b0000000000100010: out_v[37] = 10'b0001101011;
    16'b1000000000100010: out_v[37] = 10'b1100100111;
    16'b1000000000100110: out_v[37] = 10'b1001101010;
    16'b1000000000000110: out_v[37] = 10'b0110110111;
    16'b0000000000100110: out_v[37] = 10'b1011000100;
    16'b0000000000000000: out_v[37] = 10'b1101100000;
    16'b0000000000000010: out_v[37] = 10'b1101010010;
    16'b0001000000100000: out_v[37] = 10'b0010110111;
    16'b1000000000000010: out_v[37] = 10'b1011110001;
    16'b1000000000100000: out_v[37] = 10'b0011011000;
    16'b0000000000100100: out_v[37] = 10'b0011010101;
    16'b1000000000100100: out_v[37] = 10'b1101001100;
    16'b0000000000000100: out_v[37] = 10'b1100100100;
    16'b1001000000000000: out_v[37] = 10'b0000110100;
    16'b1000000000000100: out_v[37] = 10'b1111000010;
    16'b1000000000000000: out_v[37] = 10'b0010101110;
    16'b1000000000010100: out_v[37] = 10'b0111100101;
    16'b1001000000010010: out_v[37] = 10'b0010111111;
    16'b1000000000000001: out_v[37] = 10'b1010110110;
    16'b1000000000010000: out_v[37] = 10'b1000011001;
    16'b0001000000010010: out_v[37] = 10'b0000010011;
    16'b1001000000010000: out_v[37] = 10'b1111100100;
    16'b0001000000010110: out_v[37] = 10'b0000110110;
    16'b1001000000010110: out_v[37] = 10'b0101100101;
    16'b1000000000010110: out_v[37] = 10'b1010101010;
    16'b0001000000010000: out_v[37] = 10'b0010100110;
    16'b0000000000010110: out_v[37] = 10'b1010110111;
    16'b1001000000010100: out_v[37] = 10'b1010111001;
    16'b0001000000000000: out_v[37] = 10'b1110100101;
    16'b1000000000010010: out_v[37] = 10'b1010001100;
    16'b0001000000010100: out_v[37] = 10'b0100010111;
    16'b1001000000100100: out_v[37] = 10'b0001010001;
    16'b0000000000000110: out_v[37] = 10'b0010111101;
    16'b0000000000010000: out_v[37] = 10'b0000001001;
    16'b1000000000110010: out_v[37] = 10'b0110100101;
    16'b0001000000100110: out_v[37] = 10'b1110000110;
    16'b0000010010100100: out_v[37] = 10'b0100111100;
    16'b1000000000110110: out_v[37] = 10'b1010100110;
    16'b0001000000100100: out_v[37] = 10'b0110001101;
    16'b0001010010100100: out_v[37] = 10'b1001011010;
    16'b0000010010100110: out_v[37] = 10'b0110001011;
    16'b1000000000110000: out_v[37] = 10'b0110101010;
    16'b0000000010100100: out_v[37] = 10'b1001011011;
    16'b0000000000110000: out_v[37] = 10'b1101100001;
    16'b1000000000110100: out_v[37] = 10'b0111110110;
    16'b0000000010100110: out_v[37] = 10'b1101001111;
    16'b0000000010100000: out_v[37] = 10'b1010100110;
    16'b0001000010100110: out_v[37] = 10'b1001001010;
    16'b1000000010100110: out_v[37] = 10'b0011001011;
    16'b0001000000000010: out_v[37] = 10'b1001011001;
    16'b1001010010000000: out_v[37] = 10'b1001110111;
    16'b0001010010000000: out_v[37] = 10'b0110111001;
    16'b0001000010000000: out_v[37] = 10'b0101001011;
    16'b0001010010100000: out_v[37] = 10'b0001011001;
    16'b1001010010100000: out_v[37] = 10'b0111011111;
    16'b1001000010000000: out_v[37] = 10'b0100100100;
    16'b0000000010000110: out_v[37] = 10'b0000111101;
    16'b0001000000100010: out_v[37] = 10'b1110101000;
    16'b0000000010000100: out_v[37] = 10'b0110101101;
    16'b1001000000110000: out_v[37] = 10'b1111100101;
    16'b0001000000110000: out_v[37] = 10'b1010101101;
    16'b1000010010000100: out_v[37] = 10'b1001111110;
    16'b1001010010000001: out_v[37] = 10'b1001101111;
    16'b1011010010000110: out_v[37] = 10'b0111110010;
    16'b1011010010000100: out_v[37] = 10'b1011101011;
    16'b1001010010100100: out_v[37] = 10'b1001011010;
    16'b0000100000100110: out_v[37] = 10'b1011111010;
    16'b1000100000100110: out_v[37] = 10'b0111111101;
    16'b1000000000101010: out_v[37] = 10'b0100011110;
    16'b0000100000000010: out_v[37] = 10'b1001001101;
    16'b1000000000101000: out_v[37] = 10'b1101110110;
    16'b1000100000000110: out_v[37] = 10'b1101000010;
    16'b0000100000000110: out_v[37] = 10'b1100001111;
    16'b0000100000100010: out_v[37] = 10'b1001111101;
    16'b0000100000100000: out_v[37] = 10'b0011000110;
    16'b1000010010100110: out_v[37] = 10'b1100010111;
    16'b0001100000000010: out_v[37] = 10'b1001010010;
    default: out_v[37] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1000000000110000: out_v[38] = 10'b0010101011;
    16'b0000000000110000: out_v[38] = 10'b1110100000;
    16'b1000000001111000: out_v[38] = 10'b0100011101;
    16'b0000000000101000: out_v[38] = 10'b0100011111;
    16'b1000000000000000: out_v[38] = 10'b1100101100;
    16'b1000000000111000: out_v[38] = 10'b0110100111;
    16'b0000000001111000: out_v[38] = 10'b1101010011;
    16'b0000000001011000: out_v[38] = 10'b0001011011;
    16'b1000000001110000: out_v[38] = 10'b0110010000;
    16'b0000000000010000: out_v[38] = 10'b1001001010;
    16'b1000000000011000: out_v[38] = 10'b1011001001;
    16'b0000000000100000: out_v[38] = 10'b1111011001;
    16'b0000000000111000: out_v[38] = 10'b1000100001;
    16'b0000000000000000: out_v[38] = 10'b1101110010;
    16'b0000000001101000: out_v[38] = 10'b0011011001;
    16'b0000000000001000: out_v[38] = 10'b1010110100;
    16'b1000000000010000: out_v[38] = 10'b1001011011;
    16'b1000000001001000: out_v[38] = 10'b1001100000;
    16'b1000000000101000: out_v[38] = 10'b0010111000;
    16'b1000000001101000: out_v[38] = 10'b0101010111;
    16'b1000000000100000: out_v[38] = 10'b0001001011;
    16'b0000000000011000: out_v[38] = 10'b1001111011;
    16'b0000000001001000: out_v[38] = 10'b1011010011;
    16'b1000000000001000: out_v[38] = 10'b0001010110;
    16'b1000000001011000: out_v[38] = 10'b1101101010;
    16'b0000000001110000: out_v[38] = 10'b1101010111;
    16'b1010000000100000: out_v[38] = 10'b0101110111;
    16'b0000000000100010: out_v[38] = 10'b0110001010;
    16'b0000000000110010: out_v[38] = 10'b0101001001;
    16'b0010000000100000: out_v[38] = 10'b0101010111;
    16'b0010000000001000: out_v[38] = 10'b1000110010;
    16'b0010000000000000: out_v[38] = 10'b1000100111;
    16'b0010000000101000: out_v[38] = 10'b1110100010;
    16'b0010000000110000: out_v[38] = 10'b1010100001;
    16'b1000000001000000: out_v[38] = 10'b1001001111;
    16'b0000000010000000: out_v[38] = 10'b1111101011;
    16'b1000000000110010: out_v[38] = 10'b0011100000;
    16'b1000000000100010: out_v[38] = 10'b1111100011;
    16'b0010000000010000: out_v[38] = 10'b0111011010;
    16'b1000000000010010: out_v[38] = 10'b1001010111;
    16'b0010000000111000: out_v[38] = 10'b1001100111;
    default: out_v[38] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000000001001: out_v[39] = 10'b1101001000;
    16'b0000000000110111: out_v[39] = 10'b1001001001;
    16'b0000000000110101: out_v[39] = 10'b1011010110;
    16'b0000100000100100: out_v[39] = 10'b0011011110;
    16'b0000100000000000: out_v[39] = 10'b0001100100;
    16'b0000000000110001: out_v[39] = 10'b1000001111;
    16'b0000000000100101: out_v[39] = 10'b0101001001;
    16'b0000100000000100: out_v[39] = 10'b0001100111;
    16'b0000100000100000: out_v[39] = 10'b1000100010;
    16'b0000100000100101: out_v[39] = 10'b1110010111;
    16'b0000100000110001: out_v[39] = 10'b1011011110;
    16'b0000100000100111: out_v[39] = 10'b1100101011;
    16'b0000000000001100: out_v[39] = 10'b1110101111;
    16'b0000000000000100: out_v[39] = 10'b0110111001;
    16'b0000100000100110: out_v[39] = 10'b0100101001;
    16'b0000100000110100: out_v[39] = 10'b0001000100;
    16'b0000000000100100: out_v[39] = 10'b1101101010;
    16'b0000100000100001: out_v[39] = 10'b1110001101;
    16'b0000100000000001: out_v[39] = 10'b1110011011;
    16'b0000000000001101: out_v[39] = 10'b0110001011;
    16'b0000000000100111: out_v[39] = 10'b0110010101;
    16'b0000000000110011: out_v[39] = 10'b1001110100;
    16'b0000100000110000: out_v[39] = 10'b1010100110;
    16'b0000100000110101: out_v[39] = 10'b0010111101;
    16'b0000100000110110: out_v[39] = 10'b0100001111;
    16'b0000000000000111: out_v[39] = 10'b1011110001;
    16'b0000000000100110: out_v[39] = 10'b0010001011;
    16'b0000000000100000: out_v[39] = 10'b1011101011;
    16'b0000000000000001: out_v[39] = 10'b1100000101;
    16'b0000000000000101: out_v[39] = 10'b1010000101;
    16'b0000000100100101: out_v[39] = 10'b0111000011;
    16'b0000000000000000: out_v[39] = 10'b0010110110;
    16'b0000000000001000: out_v[39] = 10'b0011100111;
    16'b0000100000110111: out_v[39] = 10'b1010110100;
    16'b0000000000110100: out_v[39] = 10'b1011000110;
    16'b0000000100110101: out_v[39] = 10'b1000111001;
    16'b0001000000001100: out_v[39] = 10'b0111100011;
    16'b0000100000000101: out_v[39] = 10'b0100101100;
    16'b0000000000100001: out_v[39] = 10'b0101001100;
    16'b0000000000001111: out_v[39] = 10'b0010101111;
    16'b0000000000101101: out_v[39] = 10'b1011110101;
    16'b0000000000111001: out_v[39] = 10'b0111010011;
    16'b0000000000101001: out_v[39] = 10'b0000011011;
    16'b0000000000010001: out_v[39] = 10'b0010010110;
    16'b0000000000110000: out_v[39] = 10'b1001110110;
    16'b0000000000010000: out_v[39] = 10'b0100010111;
    16'b0000000000000010: out_v[39] = 10'b1001010011;
    16'b0000000000000011: out_v[39] = 10'b1011011010;
    16'b0000000000011001: out_v[39] = 10'b0101001001;
    16'b0001000000110001: out_v[39] = 10'b1110010100;
    16'b0000100000010000: out_v[39] = 10'b0100001001;
    16'b0000000000010101: out_v[39] = 10'b0110100110;
    16'b0000000000010100: out_v[39] = 10'b0111110010;
    16'b0000100000010001: out_v[39] = 10'b0101011010;
    16'b0000100000010100: out_v[39] = 10'b0000100101;
    16'b0001100000110000: out_v[39] = 10'b0111000110;
    16'b0000100000010110: out_v[39] = 10'b1011011110;
    16'b0000100000110010: out_v[39] = 10'b1111001100;
    16'b0001000000001001: out_v[39] = 10'b1100000110;
    16'b0001000000101001: out_v[39] = 10'b0100110101;
    16'b0000000000011000: out_v[39] = 10'b1000110011;
    16'b0001000000001000: out_v[39] = 10'b0110001011;
    16'b0000000000110010: out_v[39] = 10'b0100111100;
    16'b0000000000111000: out_v[39] = 10'b1100010000;
    16'b0001000000010100: out_v[39] = 10'b1000100111;
    16'b0000000000111010: out_v[39] = 10'b1100101010;
    16'b0001000000000100: out_v[39] = 10'b0010011011;
    16'b0001000000010001: out_v[39] = 10'b0111010001;
    16'b0001000000000000: out_v[39] = 10'b0100111101;
    16'b0000000000110110: out_v[39] = 10'b0100011010;
    16'b0000000000011100: out_v[39] = 10'b1100111101;
    16'b0001000000010000: out_v[39] = 10'b1010110010;
    16'b0001000000000001: out_v[39] = 10'b1011000011;
    16'b0000100000010101: out_v[39] = 10'b1110011010;
    16'b0000000000011101: out_v[39] = 10'b1111011110;
    16'b0000000000011110: out_v[39] = 10'b1011100110;
    16'b0000000000000110: out_v[39] = 10'b1111111000;
    16'b0000000000111100: out_v[39] = 10'b1001011000;
    16'b0000000000010110: out_v[39] = 10'b1110110010;
    16'b0000000000111101: out_v[39] = 10'b0011011010;
    16'b0000000000111110: out_v[39] = 10'b1001100111;
    16'b0000000000001010: out_v[39] = 10'b0111010010;
    16'b0000000000011011: out_v[39] = 10'b1101010110;
    16'b0000000000100010: out_v[39] = 10'b0101000110;
    16'b0000000000001011: out_v[39] = 10'b0010100101;
    16'b0000000000100011: out_v[39] = 10'b0000110111;
    16'b0000000000111011: out_v[39] = 10'b1010100011;
    16'b0000000000010011: out_v[39] = 10'b0100110110;
    16'b0000000000011010: out_v[39] = 10'b0000010001;
    16'b0000100000100010: out_v[39] = 10'b1000011111;
    16'b1000100000100000: out_v[39] = 10'b1001010110;
    16'b1000100000110000: out_v[39] = 10'b0111110000;
    16'b1000100000110100: out_v[39] = 10'b0111000100;
    16'b1000100000110001: out_v[39] = 10'b1110010011;
    16'b1000100000110101: out_v[39] = 10'b0011101110;
    16'b1000100000100001: out_v[39] = 10'b1110111011;
    16'b0000000010011001: out_v[39] = 10'b1101001000;
    16'b0000000010111001: out_v[39] = 10'b0011011011;
    16'b0000000010010001: out_v[39] = 10'b1101101111;
    16'b0000000010000001: out_v[39] = 10'b0011100000;
    16'b0000000100111001: out_v[39] = 10'b0111010111;
    16'b0000000010001001: out_v[39] = 10'b1111010101;
    16'b0000000011011001: out_v[39] = 10'b1100000101;
    16'b0000000100110001: out_v[39] = 10'b0101001111;
    16'b0000000000010010: out_v[39] = 10'b0110011011;
    16'b0001000000111001: out_v[39] = 10'b0001111111;
    16'b0000000000101000: out_v[39] = 10'b0100100101;
    16'b0001000000111000: out_v[39] = 10'b1100101110;
    16'b0000000010011000: out_v[39] = 10'b1011000101;
    16'b0001000000000101: out_v[39] = 10'b0010111000;
    16'b0001000100000101: out_v[39] = 10'b1110001111;
    16'b0001000000010101: out_v[39] = 10'b1001011111;
    default: out_v[39] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000010010001: out_v[40] = 10'b1110000101;
    16'b0000000011110011: out_v[40] = 10'b0011110010;
    16'b1000000101110011: out_v[40] = 10'b0011110011;
    16'b0000000010110001: out_v[40] = 10'b0101010110;
    16'b0000000001110010: out_v[40] = 10'b1110111011;
    16'b0000110011110011: out_v[40] = 10'b1011110001;
    16'b0000100010110001: out_v[40] = 10'b0011010001;
    16'b0000000000110001: out_v[40] = 10'b1000111001;
    16'b0000000100110001: out_v[40] = 10'b0110011011;
    16'b0000100011100011: out_v[40] = 10'b1000011111;
    16'b0000000110010001: out_v[40] = 10'b1110101101;
    16'b1000000001110011: out_v[40] = 10'b0110110111;
    16'b1000000101110000: out_v[40] = 10'b1110001010;
    16'b0000000011110010: out_v[40] = 10'b0010110010;
    16'b1100000101110011: out_v[40] = 10'b1101000110;
    16'b1000000001110001: out_v[40] = 10'b1100111100;
    16'b1000000111110001: out_v[40] = 10'b1000101100;
    16'b1100000101111001: out_v[40] = 10'b0100001011;
    16'b1100000001110011: out_v[40] = 10'b0111111010;
    16'b0000100010110011: out_v[40] = 10'b1111110010;
    16'b1000000101110001: out_v[40] = 10'b1000101101;
    16'b1000000100110001: out_v[40] = 10'b1001010111;
    16'b0000010011110011: out_v[40] = 10'b0011101010;
    16'b1000000101111001: out_v[40] = 10'b0100001101;
    16'b1100000011110011: out_v[40] = 10'b1011111110;
    16'b0000100011110011: out_v[40] = 10'b0010001101;
    16'b0001010011110011: out_v[40] = 10'b0001111101;
    16'b1100000101111011: out_v[40] = 10'b0110011010;
    16'b1000000101110010: out_v[40] = 10'b1011011110;
    16'b0000000010110011: out_v[40] = 10'b1111011011;
    16'b0000000011100011: out_v[40] = 10'b1101001110;
    16'b1000000100111001: out_v[40] = 10'b1001101011;
    16'b0000000011110001: out_v[40] = 10'b1010100110;
    16'b0000000001110011: out_v[40] = 10'b0101110111;
    16'b0000000000010001: out_v[40] = 10'b1000001110;
    16'b0000100010010001: out_v[40] = 10'b1001100011;
    16'b0000000001110001: out_v[40] = 10'b1010111110;
    16'b1100000001111001: out_v[40] = 10'b0101001111;
    16'b1100000001110001: out_v[40] = 10'b1011001110;
    16'b0000000100010001: out_v[40] = 10'b1010010101;
    16'b1100000101110001: out_v[40] = 10'b1010100111;
    16'b0000000001110000: out_v[40] = 10'b0110111010;
    16'b1000000100010001: out_v[40] = 10'b1001001101;
    16'b0000100011110001: out_v[40] = 10'b1100100110;
    16'b1000000001110010: out_v[40] = 10'b0011100111;
    16'b0000000010010000: out_v[40] = 10'b1001000111;
    16'b0000000000000000: out_v[40] = 10'b0101010011;
    16'b0000100100000000: out_v[40] = 10'b0101111010;
    16'b0000100000000000: out_v[40] = 10'b1110111001;
    16'b0000100010010000: out_v[40] = 10'b1011000000;
    16'b0000100000010000: out_v[40] = 10'b1100011111;
    16'b0000100010000000: out_v[40] = 10'b0010011111;
    16'b0000100110000000: out_v[40] = 10'b0011001111;
    16'b0001000000000001: out_v[40] = 10'b1100000111;
    16'b0000100000010001: out_v[40] = 10'b1101000000;
    16'b0000000000000001: out_v[40] = 10'b1000010100;
    16'b0000000000010000: out_v[40] = 10'b1110000100;
    16'b0000100010000001: out_v[40] = 10'b1101100001;
    16'b0000100000000001: out_v[40] = 10'b1011001011;
    16'b0000000100000000: out_v[40] = 10'b0101010111;
    16'b0000100110010000: out_v[40] = 10'b0011110110;
    16'b0000000100011001: out_v[40] = 10'b1001000110;
    16'b0100000100110011: out_v[40] = 10'b1111001011;
    16'b1100000100011001: out_v[40] = 10'b1100001101;
    16'b0000000100110011: out_v[40] = 10'b1011100110;
    16'b1000000100011001: out_v[40] = 10'b1101000110;
    16'b0000000100010000: out_v[40] = 10'b1110101001;
    16'b1100000000001000: out_v[40] = 10'b1101101101;
    16'b0000000100000001: out_v[40] = 10'b0110100101;
    16'b0100000000110011: out_v[40] = 10'b1111101111;
    16'b0000000100010011: out_v[40] = 10'b1101101001;
    16'b0000000000110011: out_v[40] = 10'b1000100111;
    16'b1000000000011001: out_v[40] = 10'b0000110011;
    16'b0100000100110001: out_v[40] = 10'b1110011011;
    16'b0100000100011001: out_v[40] = 10'b0101110111;
    16'b0000000100110010: out_v[40] = 10'b0110111001;
    16'b0000000000110010: out_v[40] = 10'b1101010001;
    16'b1100000100111001: out_v[40] = 10'b0110100011;
    16'b1100000100111011: out_v[40] = 10'b1111010011;
    16'b0000010000110011: out_v[40] = 10'b1111110110;
    16'b1000000100011011: out_v[40] = 10'b1100011011;
    16'b0000010100110010: out_v[40] = 10'b0011111011;
    16'b1000000000010001: out_v[40] = 10'b0011011101;
    16'b0100000100010001: out_v[40] = 10'b0011010011;
    16'b1000000100010000: out_v[40] = 10'b1001001100;
    16'b1100100110011001: out_v[40] = 10'b0101010100;
    16'b0000010000010011: out_v[40] = 10'b0011001101;
    16'b1000000100011000: out_v[40] = 10'b1000110111;
    16'b0000010000110010: out_v[40] = 10'b0110111011;
    16'b0000000101110010: out_v[40] = 10'b1110111001;
    16'b0000100110010001: out_v[40] = 10'b0110111000;
    16'b0000110010010011: out_v[40] = 10'b1011101100;
    16'b1000100110011001: out_v[40] = 10'b1011010100;
    16'b0000110110010011: out_v[40] = 10'b0101110001;
    16'b1000100110010011: out_v[40] = 10'b0011011111;
    16'b0000100110011001: out_v[40] = 10'b0000101111;
    16'b1000100110010001: out_v[40] = 10'b0111011000;
    16'b0000110110010001: out_v[40] = 10'b0010010001;
    16'b1001100110011001: out_v[40] = 10'b1111010111;
    16'b1000100010011001: out_v[40] = 10'b1100010000;
    16'b0000100110010011: out_v[40] = 10'b0011111011;
    16'b1000100110011000: out_v[40] = 10'b1100110001;
    16'b0000100110010010: out_v[40] = 10'b1111110001;
    16'b1000100110011011: out_v[40] = 10'b0110110011;
    16'b1000100010010001: out_v[40] = 10'b1100100011;
    16'b1000100010001000: out_v[40] = 10'b0111001011;
    16'b1000100110001000: out_v[40] = 10'b0110001101;
    16'b0000100110001000: out_v[40] = 10'b1010001010;
    16'b0000110110010010: out_v[40] = 10'b1111001110;
    16'b1000000110011001: out_v[40] = 10'b0111111011;
    16'b0000100010010011: out_v[40] = 10'b1010111000;
    16'b0000100110011000: out_v[40] = 10'b1001011110;
    16'b0000100110110001: out_v[40] = 10'b0010001110;
    16'b1000000000111001: out_v[40] = 10'b1110110000;
    16'b0000000010000000: out_v[40] = 10'b0011010000;
    16'b1000000000100001: out_v[40] = 10'b1111100010;
    16'b1000000000000001: out_v[40] = 10'b0011110001;
    16'b1000000000101001: out_v[40] = 10'b0111101000;
    16'b0000000010000001: out_v[40] = 10'b0010110101;
    16'b0000000110100000: out_v[40] = 10'b1100101001;
    16'b1000000000101000: out_v[40] = 10'b0011011111;
    16'b0000000000100001: out_v[40] = 10'b1000100100;
    16'b1000000000000000: out_v[40] = 10'b1111001100;
    16'b0000000010100000: out_v[40] = 10'b0110010011;
    16'b1000000100000000: out_v[40] = 10'b1000100010;
    16'b0000000000100000: out_v[40] = 10'b0011110110;
    16'b1000000000100000: out_v[40] = 10'b0110010010;
    16'b1000000000001001: out_v[40] = 10'b0011111011;
    16'b1000000000001000: out_v[40] = 10'b0011100101;
    16'b0000000011100000: out_v[40] = 10'b1110110100;
    16'b0000000001100000: out_v[40] = 10'b0001011100;
    16'b1000000001101000: out_v[40] = 10'b0100110011;
    16'b0000000010100001: out_v[40] = 10'b1110101100;
    16'b0000100010100000: out_v[40] = 10'b0110101110;
    16'b0000100010100001: out_v[40] = 10'b0001110011;
    16'b0000000100100000: out_v[40] = 10'b0010110101;
    16'b0000000110000001: out_v[40] = 10'b0000110101;
    16'b1000000100100000: out_v[40] = 10'b0111011100;
    16'b1000000101100000: out_v[40] = 10'b0001010110;
    16'b0000000110000000: out_v[40] = 10'b0011111011;
    16'b1000000000110001: out_v[40] = 10'b1101001000;
    16'b0000000010110000: out_v[40] = 10'b0011010111;
    16'b1000000001100000: out_v[40] = 10'b0110010011;
    16'b0000100010000010: out_v[40] = 10'b0000011101;
    16'b0000000010000011: out_v[40] = 10'b1101011110;
    16'b1000000110010001: out_v[40] = 10'b1000110100;
    16'b0000000000000011: out_v[40] = 10'b1111101001;
    16'b0000100010010010: out_v[40] = 10'b1100101111;
    16'b1000100110010000: out_v[40] = 10'b0110100000;
    16'b0000100010000011: out_v[40] = 10'b1111110100;
    16'b0000000010010011: out_v[40] = 10'b0111111111;
    16'b1000100010010000: out_v[40] = 10'b0000111000;
    16'b1000000110010000: out_v[40] = 10'b1010101011;
    16'b1000000010010000: out_v[40] = 10'b1100101010;
    16'b0000000110010000: out_v[40] = 10'b1001101000;
    16'b1000000000010000: out_v[40] = 10'b1010111000;
    16'b1000000010010001: out_v[40] = 10'b0010001111;
    16'b1000000110011000: out_v[40] = 10'b0011110011;
    16'b1000000101000000: out_v[40] = 10'b1111101010;
    16'b1100000001101000: out_v[40] = 10'b0010010111;
    16'b1100000100100000: out_v[40] = 10'b1111001001;
    16'b1000000110000000: out_v[40] = 10'b0111010111;
    16'b0000000000110000: out_v[40] = 10'b1001000101;
    16'b1100000101100000: out_v[40] = 10'b0111111011;
    16'b1100000101101000: out_v[40] = 10'b1111011100;
    16'b0000000011110000: out_v[40] = 10'b1011111000;
    16'b0000000101000000: out_v[40] = 10'b0001011010;
    16'b0000100010110000: out_v[40] = 10'b0101110010;
    16'b1000000101101000: out_v[40] = 10'b0010011111;
    16'b1000000010000001: out_v[40] = 10'b0011101010;
    16'b1000000001001001: out_v[40] = 10'b0010101011;
    16'b1000000001000001: out_v[40] = 10'b1001101011;
    16'b1001000000000001: out_v[40] = 10'b1111111111;
    16'b1000100010000001: out_v[40] = 10'b1000110100;
    16'b0001000000010001: out_v[40] = 10'b0111111000;
    16'b1000000001100001: out_v[40] = 10'b1101110111;
    default: out_v[40] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1110000110010000: out_v[41] = 10'b0000011111;
    16'b1110000010011100: out_v[41] = 10'b0111010010;
    16'b1010000110001000: out_v[41] = 10'b0001111001;
    16'b0110000100010000: out_v[41] = 10'b1101110000;
    16'b1110000010010000: out_v[41] = 10'b1101001011;
    16'b1010000110100000: out_v[41] = 10'b1010000111;
    16'b1110000011011000: out_v[41] = 10'b0000011101;
    16'b1010000010000000: out_v[41] = 10'b0101010010;
    16'b0010000100001000: out_v[41] = 10'b0111000110;
    16'b0110000110010000: out_v[41] = 10'b0101110110;
    16'b1100000010010100: out_v[41] = 10'b1001100111;
    16'b1010000011001000: out_v[41] = 10'b1011110010;
    16'b1110000010011000: out_v[41] = 10'b0100100000;
    16'b1010000010001000: out_v[41] = 10'b0010100011;
    16'b0010000110001000: out_v[41] = 10'b0100010100;
    16'b0010000110000000: out_v[41] = 10'b0000111111;
    16'b1110000111010000: out_v[41] = 10'b1100001000;
    16'b0010000100000000: out_v[41] = 10'b1101001011;
    16'b1010000110000000: out_v[41] = 10'b1010011111;
    16'b1110000010010100: out_v[41] = 10'b0000100101;
    16'b0010000000000000: out_v[41] = 10'b1001011011;
    16'b1000000010001100: out_v[41] = 10'b0011100001;
    16'b1000000011001100: out_v[41] = 10'b1101110011;
    16'b0010000110100000: out_v[41] = 10'b1110001011;
    16'b0010000110101000: out_v[41] = 10'b1000110101;
    16'b1010000110101000: out_v[41] = 10'b0011010011;
    16'b1110000011011100: out_v[41] = 10'b1001110000;
    16'b1110000110011000: out_v[41] = 10'b1100110011;
    16'b1010000111000000: out_v[41] = 10'b1110111110;
    16'b1010000111001000: out_v[41] = 10'b1101100010;
    16'b1100000010010000: out_v[41] = 10'b1000010010;
    16'b0110000010010000: out_v[41] = 10'b1100100001;
    16'b1010000011000000: out_v[41] = 10'b0001111001;
    16'b1110000011010000: out_v[41] = 10'b0011010110;
    16'b0100000100010000: out_v[41] = 10'b0001110011;
    16'b1100000110010000: out_v[41] = 10'b1110001001;
    16'b0010000100100000: out_v[41] = 10'b1111101101;
    16'b1010000010001100: out_v[41] = 10'b1011000011;
    16'b1010000110001100: out_v[41] = 10'b1101001110;
    16'b1000000110001100: out_v[41] = 10'b1011110011;
    16'b1010000011001100: out_v[41] = 10'b1010110011;
    16'b0010000010000000: out_v[41] = 10'b0100011101;
    16'b0110000000010000: out_v[41] = 10'b0110000111;
    16'b0000000000000000: out_v[41] = 10'b0110010010;
    16'b1000000010000000: out_v[41] = 10'b1010011110;
    16'b0010000000000100: out_v[41] = 10'b1100010011;
    16'b1000000110000000: out_v[41] = 10'b1110001000;
    16'b0000000100000000: out_v[41] = 10'b0100110000;
    16'b1010000000000000: out_v[41] = 10'b0111001000;
    16'b1000000000000000: out_v[41] = 10'b1111100110;
    16'b0000000010000000: out_v[41] = 10'b1101010001;
    16'b0000000110000000: out_v[41] = 10'b0110101100;
    16'b0010000000100000: out_v[41] = 10'b1110001110;
    16'b0100000000010000: out_v[41] = 10'b0010011001;
    16'b1000000110100000: out_v[41] = 10'b1010110101;
    16'b0110000001010000: out_v[41] = 10'b0101010100;
    16'b0110000100010100: out_v[41] = 10'b1111110000;
    16'b0110000110010100: out_v[41] = 10'b1111100100;
    16'b0110000101010000: out_v[41] = 10'b0001110101;
    16'b0110000111010000: out_v[41] = 10'b1010111010;
    16'b0010000100000100: out_v[41] = 10'b1110110100;
    16'b0110000000110000: out_v[41] = 10'b1001100110;
    16'b0110000110110000: out_v[41] = 10'b0101110110;
    16'b0110000100110000: out_v[41] = 10'b0101110110;
    16'b1110000110010100: out_v[41] = 10'b1011011011;
    16'b0010000110000100: out_v[41] = 10'b0011110100;
    16'b0110000011010000: out_v[41] = 10'b1010101010;
    16'b1010000010100000: out_v[41] = 10'b1000110110;
    16'b1110000110110000: out_v[41] = 10'b1100010110;
    16'b0100000100010100: out_v[41] = 10'b1111010011;
    16'b0100000110010100: out_v[41] = 10'b0101001010;
    16'b0100000110010000: out_v[41] = 10'b1100110100;
    16'b0000000100000100: out_v[41] = 10'b0101010100;
    16'b0100000101010100: out_v[41] = 10'b1010101000;
    16'b1000000110000100: out_v[41] = 10'b1000001011;
    16'b0000000000000100: out_v[41] = 10'b0000011010;
    16'b0000000110000100: out_v[41] = 10'b0010110111;
    16'b1110000000010000: out_v[41] = 10'b1011001001;
    16'b0100000111010100: out_v[41] = 10'b0111111110;
    16'b1100000110010100: out_v[41] = 10'b0101011001;
    16'b0100000000010100: out_v[41] = 10'b0011011010;
    16'b0010000001000000: out_v[41] = 10'b1110011011;
    16'b1110000100010000: out_v[41] = 10'b0100110010;
    16'b0100000110011000: out_v[41] = 10'b1010000110;
    16'b0100000100011000: out_v[41] = 10'b0000011000;
    16'b0100000010010000: out_v[41] = 10'b1000110011;
    16'b1100000010011000: out_v[41] = 10'b1000010000;
    16'b0100000000011000: out_v[41] = 10'b1010001111;
    16'b0010000000001000: out_v[41] = 10'b1001101000;
    16'b1000000110001000: out_v[41] = 10'b0001100100;
    16'b1010000000001000: out_v[41] = 10'b1001110001;
    16'b1000000010000100: out_v[41] = 10'b1010100010;
    16'b1010000010000100: out_v[41] = 10'b0110110000;
    16'b1000000010001000: out_v[41] = 10'b0000100111;
    16'b0000000000001000: out_v[41] = 10'b0010100000;
    16'b1110001010010000: out_v[41] = 10'b0011101110;
    16'b1110001110010000: out_v[41] = 10'b0110110111;
    16'b0100000100110000: out_v[41] = 10'b0111100011;
    16'b0110001100010000: out_v[41] = 10'b1001111010;
    16'b1010001010000000: out_v[41] = 10'b0101100011;
    16'b1000001010000000: out_v[41] = 10'b1111000101;
    16'b0110001010010000: out_v[41] = 10'b1001011111;
    16'b0110001110010000: out_v[41] = 10'b0111111010;
    16'b1100000000010000: out_v[41] = 10'b1000001010;
    16'b1110000110011100: out_v[41] = 10'b0011001110;
    16'b1100000000011000: out_v[41] = 10'b1000011010;
    16'b1100000110011000: out_v[41] = 10'b0111101010;
    16'b1100000010011100: out_v[41] = 10'b0101011011;
    16'b0110000110011000: out_v[41] = 10'b0111010010;
    16'b0110000110011100: out_v[41] = 10'b0110011001;
    16'b0110000100011000: out_v[41] = 10'b1101010000;
    default: out_v[41] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000011100000001: out_v[42] = 10'b0111001011;
    16'b0000001100000001: out_v[42] = 10'b1000100110;
    16'b1010011100100001: out_v[42] = 10'b0100010000;
    16'b1000011100100011: out_v[42] = 10'b1011011010;
    16'b1000011100100001: out_v[42] = 10'b0001000011;
    16'b1000010100100001: out_v[42] = 10'b1101011001;
    16'b1000001100100001: out_v[42] = 10'b0011111011;
    16'b0010011100000000: out_v[42] = 10'b0010100111;
    16'b0010011100000001: out_v[42] = 10'b0100101011;
    16'b1010011100100000: out_v[42] = 10'b0010110110;
    16'b1000011100000001: out_v[42] = 10'b1000110010;
    16'b1010011000100000: out_v[42] = 10'b1101001011;
    16'b0000010100000001: out_v[42] = 10'b1001110000;
    16'b0010001100000001: out_v[42] = 10'b0010011110;
    16'b1000001100000001: out_v[42] = 10'b1010110011;
    16'b1010011100100011: out_v[42] = 10'b0011000011;
    16'b1000010100000001: out_v[42] = 10'b0101100011;
    16'b0000011000000001: out_v[42] = 10'b0110100001;
    16'b1010011000100010: out_v[42] = 10'b1001101111;
    16'b0010011000000000: out_v[42] = 10'b0000001110;
    16'b1010001000100000: out_v[42] = 10'b0001101111;
    16'b0000001000000001: out_v[42] = 10'b1011100000;
    16'b0000011100000000: out_v[42] = 10'b0111001010;
    16'b1010011000100011: out_v[42] = 10'b1001010110;
    16'b0000001000000000: out_v[42] = 10'b0001011011;
    16'b0010001100000000: out_v[42] = 10'b1101010010;
    16'b0000001100000000: out_v[42] = 10'b0111110001;
    16'b0010011100000011: out_v[42] = 10'b0001110100;
    16'b0000010000000000: out_v[42] = 10'b0011010011;
    16'b0000000000000000: out_v[42] = 10'b0100010011;
    16'b0010000000000001: out_v[42] = 10'b0011101011;
    16'b0000011000000000: out_v[42] = 10'b0001011100;
    16'b0000000000000001: out_v[42] = 10'b0010110001;
    16'b0010001000000001: out_v[42] = 10'b0000101010;
    16'b0010011000000010: out_v[42] = 10'b0001010110;
    16'b1010010000000010: out_v[42] = 10'b1010011010;
    16'b0010001000000000: out_v[42] = 10'b0010001101;
    16'b0000010000000001: out_v[42] = 10'b0011011100;
    16'b0000000000000011: out_v[42] = 10'b1101010100;
    16'b0010010000000000: out_v[42] = 10'b0000000101;
    16'b1000010000100000: out_v[42] = 10'b0100001100;
    16'b0010010000000010: out_v[42] = 10'b1011010011;
    16'b0010010000000001: out_v[42] = 10'b1100110101;
    16'b1000010000000001: out_v[42] = 10'b0010001110;
    16'b1000010000000000: out_v[42] = 10'b1010110101;
    16'b1010010000000000: out_v[42] = 10'b1000100101;
    16'b0010011000000011: out_v[42] = 10'b0000110101;
    16'b0000010000000010: out_v[42] = 10'b0100111101;
    16'b0010000000000000: out_v[42] = 10'b1011001001;
    16'b1010010000100010: out_v[42] = 10'b1101111110;
    16'b0010011000000001: out_v[42] = 10'b1100010111;
    16'b0000010000000011: out_v[42] = 10'b0010101111;
    16'b1010010000000001: out_v[42] = 10'b1010011111;
    16'b1000010000000010: out_v[42] = 10'b1101100101;
    16'b1000000000000000: out_v[42] = 10'b0000110101;
    16'b0010010000000011: out_v[42] = 10'b1100110111;
    16'b0010001000000010: out_v[42] = 10'b0000111101;
    16'b1010010000100000: out_v[42] = 10'b1011100010;
    16'b0010011010000000: out_v[42] = 10'b1001001110;
    16'b1000010000000011: out_v[42] = 10'b0011101010;
    16'b1000000000000001: out_v[42] = 10'b1101000100;
    16'b0010000000000010: out_v[42] = 10'b1101010111;
    16'b1000010000100001: out_v[42] = 10'b1110000110;
    16'b1010011000000000: out_v[42] = 10'b0011011111;
    16'b1000000000100000: out_v[42] = 10'b0111110111;
    16'b0010001010000000: out_v[42] = 10'b1001101110;
    16'b1010001100000000: out_v[42] = 10'b1111100010;
    16'b1000011000000001: out_v[42] = 10'b0110111100;
    16'b1000011000000000: out_v[42] = 10'b0010111011;
    16'b1010011100000000: out_v[42] = 10'b1001110011;
    16'b1010001000000000: out_v[42] = 10'b1010011110;
    16'b1000001000000000: out_v[42] = 10'b1110110111;
    16'b0010001000001000: out_v[42] = 10'b0011111110;
    16'b1000001000000001: out_v[42] = 10'b1111101110;
    16'b0000000100000000: out_v[42] = 10'b1010110001;
    16'b0010000100100000: out_v[42] = 10'b0100110111;
    16'b0000000100000001: out_v[42] = 10'b1100110111;
    16'b0010000000100000: out_v[42] = 10'b1011001101;
    16'b0000010100000000: out_v[42] = 10'b1100000111;
    16'b0010000100000000: out_v[42] = 10'b0100110000;
    16'b0000001100100001: out_v[42] = 10'b0111110010;
    16'b0010001100100000: out_v[42] = 10'b1101111011;
    16'b1000000100100000: out_v[42] = 10'b0011001010;
    16'b1000000100000001: out_v[42] = 10'b1101011000;
    16'b0010000100000001: out_v[42] = 10'b1010101010;
    16'b0000000010100000: out_v[42] = 10'b0111110010;
    16'b0000000100100001: out_v[42] = 10'b0000011100;
    16'b1000000100100001: out_v[42] = 10'b1111000011;
    16'b0000000000100000: out_v[42] = 10'b0101110000;
    16'b0000001100100000: out_v[42] = 10'b0011011010;
    16'b0000000100100000: out_v[42] = 10'b0010010101;
    16'b0000010100100001: out_v[42] = 10'b0010101111;
    16'b0000001000100000: out_v[42] = 10'b1100101010;
    16'b0010011100000010: out_v[42] = 10'b1110100001;
    16'b0010001100000010: out_v[42] = 10'b0111101011;
    16'b1000010100000000: out_v[42] = 10'b1101100100;
    16'b0010010100000010: out_v[42] = 10'b1111110111;
    16'b0010000100000010: out_v[42] = 10'b0111100110;
    16'b0010010100000001: out_v[42] = 10'b0010011101;
    16'b0010010100000000: out_v[42] = 10'b0100010000;
    16'b0000000011000001: out_v[42] = 10'b0111010011;
    16'b0000001011000001: out_v[42] = 10'b1001011011;
    16'b0000000001000001: out_v[42] = 10'b0111101001;
    16'b0000001001000001: out_v[42] = 10'b0011100101;
    16'b0000001101000001: out_v[42] = 10'b0011010110;
    16'b0000001010000001: out_v[42] = 10'b0011010000;
    16'b0000000101000001: out_v[42] = 10'b1100001110;
    16'b0000010000001001: out_v[42] = 10'b1011010011;
    16'b0001000101000001: out_v[42] = 10'b1100011111;
    16'b0000000010000001: out_v[42] = 10'b1111110000;
    16'b0001000001000001: out_v[42] = 10'b1011111011;
    16'b0001000011000001: out_v[42] = 10'b1001110101;
    16'b0000000000100001: out_v[42] = 10'b1111000111;
    16'b0000000101000000: out_v[42] = 10'b1000101101;
    default: out_v[42] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000000000000: out_v[43] = 10'b1111100110;
    16'b0101000100000000: out_v[43] = 10'b0111001011;
    16'b0101000100100000: out_v[43] = 10'b1011000001;
    16'b0001000100100000: out_v[43] = 10'b0100010100;
    16'b0001000000000000: out_v[43] = 10'b0100110100;
    16'b0001000100000000: out_v[43] = 10'b0100010100;
    16'b0100000100100000: out_v[43] = 10'b0110010111;
    16'b0100000000100000: out_v[43] = 10'b1101100011;
    16'b0100000000000000: out_v[43] = 10'b1100011110;
    16'b0000000100000000: out_v[43] = 10'b1011110000;
    16'b0100000100000000: out_v[43] = 10'b1000011111;
    16'b0101000000000000: out_v[43] = 10'b1110100010;
    16'b0101000000100000: out_v[43] = 10'b0010011001;
    16'b0001000000100000: out_v[43] = 10'b1010011001;
    16'b0000000100100000: out_v[43] = 10'b0011110000;
    16'b0100000001000000: out_v[43] = 10'b0000001101;
    16'b0000000101000000: out_v[43] = 10'b0011000100;
    16'b0001000001000000: out_v[43] = 10'b1000111110;
    16'b0001000101000000: out_v[43] = 10'b0011101111;
    16'b1001000100100000: out_v[43] = 10'b0100100111;
    16'b0100000101000000: out_v[43] = 10'b0110010110;
    16'b0001010000000000: out_v[43] = 10'b0000111111;
    16'b0001000101100000: out_v[43] = 10'b0110110111;
    16'b1001000100000000: out_v[43] = 10'b1111000101;
    16'b1001000000000000: out_v[43] = 10'b0011111010;
    16'b1101000000000000: out_v[43] = 10'b0001001110;
    16'b0000000001000000: out_v[43] = 10'b0111000010;
    16'b1001010000000000: out_v[43] = 10'b0111001000;
    16'b0101010000000000: out_v[43] = 10'b0010101000;
    16'b0100010000000000: out_v[43] = 10'b1111001011;
    16'b1101010000000000: out_v[43] = 10'b1101011110;
    16'b0000000101100000: out_v[43] = 10'b1011100110;
    16'b0100000000000001: out_v[43] = 10'b0111111010;
    16'b0000000100000001: out_v[43] = 10'b1101101011;
    16'b0100000100000001: out_v[43] = 10'b0111101011;
    16'b0000000000000001: out_v[43] = 10'b1111101110;
    16'b0100000010000000: out_v[43] = 10'b0010011011;
    16'b0100000110000000: out_v[43] = 10'b1011001101;
    16'b0100000110100000: out_v[43] = 10'b1001100100;
    default: out_v[43] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1010000000010000: out_v[44] = 10'b0111111101;
    16'b1000000000000001: out_v[44] = 10'b0011011101;
    16'b1000000001001001: out_v[44] = 10'b1010000011;
    16'b1010000000011001: out_v[44] = 10'b1010010111;
    16'b0000000000000000: out_v[44] = 10'b0010110000;
    16'b1000000001000001: out_v[44] = 10'b0100110001;
    16'b0010000001001001: out_v[44] = 10'b1010110110;
    16'b1010000000010001: out_v[44] = 10'b1111000000;
    16'b0000000000000001: out_v[44] = 10'b0010101110;
    16'b1000000000010011: out_v[44] = 10'b1000100011;
    16'b0000100000000001: out_v[44] = 10'b0100010100;
    16'b1010000001001000: out_v[44] = 10'b0001011101;
    16'b0010000000001000: out_v[44] = 10'b0011001101;
    16'b1010000000011000: out_v[44] = 10'b0111000011;
    16'b1010000000000001: out_v[44] = 10'b1000010101;
    16'b1000000001001000: out_v[44] = 10'b1000110010;
    16'b1010000001001001: out_v[44] = 10'b1110011000;
    16'b1000000000000000: out_v[44] = 10'b1011100011;
    16'b1000000000010001: out_v[44] = 10'b0010001111;
    16'b1010000001011001: out_v[44] = 10'b0001011011;
    16'b0000000001001001: out_v[44] = 10'b1001100110;
    16'b1010000000001001: out_v[44] = 10'b0000011110;
    16'b1001000000000001: out_v[44] = 10'b0101000011;
    16'b0010000001001000: out_v[44] = 10'b1001100011;
    16'b1000000000001001: out_v[44] = 10'b1101011011;
    16'b0000000000010000: out_v[44] = 10'b1001011011;
    16'b1000100000000001: out_v[44] = 10'b1111101011;
    16'b1000000000010000: out_v[44] = 10'b1000010011;
    16'b1010000000000000: out_v[44] = 10'b0011000011;
    16'b1000000000011001: out_v[44] = 10'b0110011011;
    16'b0000000001000001: out_v[44] = 10'b0010011011;
    16'b0001000000000001: out_v[44] = 10'b1001110101;
    16'b0000000000010001: out_v[44] = 10'b1101000100;
    16'b1000000000001000: out_v[44] = 10'b1111100011;
    16'b0010000000000000: out_v[44] = 10'b1011001110;
    16'b1010000000001000: out_v[44] = 10'b0011101011;
    16'b1000000001011001: out_v[44] = 10'b0101001101;
    16'b1000000000000011: out_v[44] = 10'b1001110010;
    16'b0000000000000010: out_v[44] = 10'b1100000010;
    16'b0000000000000011: out_v[44] = 10'b1101001010;
    16'b0010000000000010: out_v[44] = 10'b0011011101;
    16'b0010000000000011: out_v[44] = 10'b0100100010;
    16'b1000000000000010: out_v[44] = 10'b1100011101;
    16'b0000000000010011: out_v[44] = 10'b1011000000;
    16'b1000000000010010: out_v[44] = 10'b1100111100;
    16'b0010000000001010: out_v[44] = 10'b1001010010;
    16'b0010000000001011: out_v[44] = 10'b0100100000;
    16'b1000000000011011: out_v[44] = 10'b0011110110;
    16'b0000000000001001: out_v[44] = 10'b1100100011;
    16'b1000000000001011: out_v[44] = 10'b0011010000;
    16'b0000000000011011: out_v[44] = 10'b0100010100;
    16'b0000000001001011: out_v[44] = 10'b1011000010;
    16'b0000000000001011: out_v[44] = 10'b0110010100;
    16'b0000000000010010: out_v[44] = 10'b0100100111;
    16'b0000000000011001: out_v[44] = 10'b1101101110;
    16'b1001000000010011: out_v[44] = 10'b0110100111;
    16'b1000000000011010: out_v[44] = 10'b0111010110;
    16'b0010000000011011: out_v[44] = 10'b0001101111;
    16'b1000000001011011: out_v[44] = 10'b1011101100;
    16'b0000000000011010: out_v[44] = 10'b1010101000;
    16'b0001000000010011: out_v[44] = 10'b1111101110;
    16'b1000000001001011: out_v[44] = 10'b1101110110;
    16'b0000000001011011: out_v[44] = 10'b0001001000;
    16'b1010000000001011: out_v[44] = 10'b0000101011;
    16'b1001000000011011: out_v[44] = 10'b0101010111;
    16'b1010000000011011: out_v[44] = 10'b0110110010;
    16'b1001000000010001: out_v[44] = 10'b1111010100;
    16'b0000000000011110: out_v[44] = 10'b1101001111;
    16'b1001000000010010: out_v[44] = 10'b0001011110;
    16'b0000000000011111: out_v[44] = 10'b0000010110;
    16'b0001000000011011: out_v[44] = 10'b1111010011;
    16'b1001000000001011: out_v[44] = 10'b0101011101;
    16'b1010000001001011: out_v[44] = 10'b0000100111;
    16'b1010000000011010: out_v[44] = 10'b1111000100;
    16'b0010000000011010: out_v[44] = 10'b0010111000;
    16'b1001000000000011: out_v[44] = 10'b0000001011;
    16'b1001000000000000: out_v[44] = 10'b1111000011;
    16'b1010000000001010: out_v[44] = 10'b1111001000;
    16'b0000000000001000: out_v[44] = 10'b0011001010;
    16'b1001000000001001: out_v[44] = 10'b1111011010;
    16'b0010000000001001: out_v[44] = 10'b1001111101;
    16'b0000000000001010: out_v[44] = 10'b1101001011;
    16'b1011000000001010: out_v[44] = 10'b0111100011;
    16'b1011000000001000: out_v[44] = 10'b1100111010;
    16'b1001000000001000: out_v[44] = 10'b0101010011;
    16'b0010000001001010: out_v[44] = 10'b1001001111;
    16'b1001000000001010: out_v[44] = 10'b0111110111;
    16'b1010000001001010: out_v[44] = 10'b1101011011;
    16'b1000000000001010: out_v[44] = 10'b0000011111;
    16'b1010000000000010: out_v[44] = 10'b1000011111;
    16'b0010000000000001: out_v[44] = 10'b1001001100;
    16'b1010000001011010: out_v[44] = 10'b1100011000;
    16'b0000000001011010: out_v[44] = 10'b1100000000;
    16'b0010000001011010: out_v[44] = 10'b1100111010;
    16'b0000100000010011: out_v[44] = 10'b0100110001;
    16'b1000000001011010: out_v[44] = 10'b0001111000;
    16'b0010000000010010: out_v[44] = 10'b1000101010;
    16'b1010000000010010: out_v[44] = 10'b1000111110;
    16'b0010000001000010: out_v[44] = 10'b0111111011;
    16'b0010000001010010: out_v[44] = 10'b0110110011;
    16'b1010000001011000: out_v[44] = 10'b0110010111;
    16'b1000100000010011: out_v[44] = 10'b1101101001;
    16'b0000000001010010: out_v[44] = 10'b1000100110;
    16'b0010000000011000: out_v[44] = 10'b0110110011;
    16'b1000000001010010: out_v[44] = 10'b1011111000;
    16'b1010000001010010: out_v[44] = 10'b1001001110;
    16'b0010000000010000: out_v[44] = 10'b0011011000;
    16'b1000100000000011: out_v[44] = 10'b0010110011;
    16'b0010100000000010: out_v[44] = 10'b1101001111;
    16'b0010000001001011: out_v[44] = 10'b0000001111;
    16'b0000100000000011: out_v[44] = 10'b1010101111;
    16'b0010100001001010: out_v[44] = 10'b1111110000;
    16'b1000100000000010: out_v[44] = 10'b1001110111;
    16'b1000100000010001: out_v[44] = 10'b1101101110;
    16'b0000000001011111: out_v[44] = 10'b1110100101;
    16'b0000000001011001: out_v[44] = 10'b1101000010;
    16'b0010000000010011: out_v[44] = 10'b1011010101;
    16'b1010000001000000: out_v[44] = 10'b0011001000;
    16'b1000000001000000: out_v[44] = 10'b0111100001;
    16'b0000000001001000: out_v[44] = 10'b1001110011;
    16'b0000000001000000: out_v[44] = 10'b0111001010;
    16'b1000000001000011: out_v[44] = 10'b1011001001;
    16'b0010000001000000: out_v[44] = 10'b0111010101;
    16'b1010000000000011: out_v[44] = 10'b0100000001;
    16'b1010000000010011: out_v[44] = 10'b1001001010;
    16'b1010000001011011: out_v[44] = 10'b1110010011;
    16'b0010000001011011: out_v[44] = 10'b0110100110;
    16'b1000100000010010: out_v[44] = 10'b0011010111;
    16'b1000000001010011: out_v[44] = 10'b0111011110;
    16'b1000000001001010: out_v[44] = 10'b0011100110;
    16'b1000000001011000: out_v[44] = 10'b1100000110;
    16'b0000000001001010: out_v[44] = 10'b1101001111;
    16'b0010000001011000: out_v[44] = 10'b1100110010;
    16'b0000000001011000: out_v[44] = 10'b0010111010;
    default: out_v[44] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0011000000110000: out_v[45] = 10'b1110001111;
    16'b0011000000111010: out_v[45] = 10'b0110110111;
    16'b0011000010111010: out_v[45] = 10'b0101101001;
    16'b0011000010110000: out_v[45] = 10'b0001100011;
    16'b0011000000111001: out_v[45] = 10'b1000001001;
    16'b0011000000111011: out_v[45] = 10'b1001001011;
    16'b0001000000111000: out_v[45] = 10'b0001011001;
    16'b0001000000101010: out_v[45] = 10'b0111011011;
    16'b0001000010110000: out_v[45] = 10'b0111110111;
    16'b0011000000101010: out_v[45] = 10'b1111001100;
    16'b0011000010110010: out_v[45] = 10'b0100110001;
    16'b0011000000100010: out_v[45] = 10'b0010101001;
    16'b0011000000111000: out_v[45] = 10'b0000110110;
    16'b0011000010111000: out_v[45] = 10'b0011100011;
    16'b0010000010010000: out_v[45] = 10'b1011100101;
    16'b0011000000010010: out_v[45] = 10'b0010011111;
    16'b0010000010011010: out_v[45] = 10'b0101101000;
    16'b0010000010010010: out_v[45] = 10'b1110111011;
    16'b0000000010011010: out_v[45] = 10'b1000110111;
    16'b0011000000010000: out_v[45] = 10'b1010100001;
    16'b0011000000011000: out_v[45] = 10'b1100111011;
    16'b0011000000011010: out_v[45] = 10'b0011110100;
    16'b0011000000110010: out_v[45] = 10'b1001001001;
    16'b0000000010010010: out_v[45] = 10'b1000011101;
    16'b0001000000100010: out_v[45] = 10'b1011010011;
    16'b0010000000011010: out_v[45] = 10'b0100011010;
    16'b0000000010011000: out_v[45] = 10'b0010001101;
    16'b0001000000111010: out_v[45] = 10'b1000000110;
    16'b0001000010110010: out_v[45] = 10'b0110000010;
    16'b0011000000011011: out_v[45] = 10'b1010011101;
    16'b0011000000011001: out_v[45] = 10'b1000111011;
    16'b0011000010101000: out_v[45] = 10'b0011010001;
    16'b0011000010111011: out_v[45] = 10'b1101000110;
    16'b0011000010111001: out_v[45] = 10'b0011010101;
    16'b0001000000110010: out_v[45] = 10'b0011011111;
    16'b0010000010011000: out_v[45] = 10'b1110101011;
    16'b0010000010110000: out_v[45] = 10'b0111110110;
    16'b0001000010111010: out_v[45] = 10'b1111010101;
    16'b0001000010111000: out_v[45] = 10'b0001111111;
    16'b0000000010010000: out_v[45] = 10'b1001010111;
    16'b0010000000011011: out_v[45] = 10'b0101011101;
    16'b0000000000010011: out_v[45] = 10'b1011000011;
    16'b0000000000011001: out_v[45] = 10'b0010100110;
    16'b0000000000001000: out_v[45] = 10'b1001010110;
    16'b0000000000000000: out_v[45] = 10'b1100000100;
    16'b0000000000001001: out_v[45] = 10'b1001100101;
    16'b0000000000000001: out_v[45] = 10'b0101011100;
    16'b0000000000010010: out_v[45] = 10'b1011101011;
    16'b0000000000011011: out_v[45] = 10'b0001011010;
    16'b0000000000010000: out_v[45] = 10'b1011100000;
    16'b0000000000011000: out_v[45] = 10'b0101111101;
    16'b0000000010000001: out_v[45] = 10'b0111001010;
    16'b0000000000011010: out_v[45] = 10'b1110110101;
    16'b0000000000000010: out_v[45] = 10'b1111100010;
    16'b0000000010001001: out_v[45] = 10'b0101101100;
    16'b0001000000001001: out_v[45] = 10'b1010101000;
    16'b0000000000001011: out_v[45] = 10'b0111010011;
    16'b0010000010011011: out_v[45] = 10'b1000011000;
    16'b0000000010001011: out_v[45] = 10'b1101010111;
    16'b0000000000010001: out_v[45] = 10'b0000111100;
    16'b0000000010001000: out_v[45] = 10'b0010111101;
    16'b0010000010001001: out_v[45] = 10'b0111100110;
    16'b0010000000010001: out_v[45] = 10'b1100000110;
    16'b0000000010011011: out_v[45] = 10'b1000011011;
    16'b0000000010011001: out_v[45] = 10'b0110101100;
    16'b0010000000011001: out_v[45] = 10'b0110010101;
    16'b0010000010010001: out_v[45] = 10'b1001001101;
    16'b0000000000001010: out_v[45] = 10'b0011100101;
    16'b0000000010010001: out_v[45] = 10'b0101001010;
    16'b0011000010011011: out_v[45] = 10'b0000101110;
    16'b0010000000001011: out_v[45] = 10'b1110101000;
    16'b0010000010011001: out_v[45] = 10'b0010100111;
    16'b0010000000010011: out_v[45] = 10'b1110000010;
    16'b0010000000000001: out_v[45] = 10'b0100010100;
    16'b0001000010011011: out_v[45] = 10'b1011001001;
    16'b0010000010010011: out_v[45] = 10'b0111101111;
    16'b0000000010010011: out_v[45] = 10'b0001111110;
    16'b0100000010001001: out_v[45] = 10'b1110101101;
    16'b0000000000000011: out_v[45] = 10'b0000101001;
    16'b0001000000011011: out_v[45] = 10'b1010100111;
    16'b0000000010000000: out_v[45] = 10'b0011011101;
    16'b0000000010001010: out_v[45] = 10'b1011010101;
    16'b0010000010001011: out_v[45] = 10'b0001111110;
    16'b0000000010000010: out_v[45] = 10'b1010001101;
    16'b0010000010000010: out_v[45] = 10'b1011001110;
    16'b0000000010000011: out_v[45] = 10'b1111010111;
    16'b0010000010000000: out_v[45] = 10'b1010001101;
    16'b0011000000110001: out_v[45] = 10'b0100000011;
    16'b0001000010100001: out_v[45] = 10'b0111110010;
    16'b0001000000101001: out_v[45] = 10'b0010011110;
    16'b0011000000101001: out_v[45] = 10'b0011110010;
    16'b0000000010110001: out_v[45] = 10'b0111000010;
    16'b0000000000110001: out_v[45] = 10'b0111000101;
    16'b0001000000111001: out_v[45] = 10'b0110000101;
    16'b0001000000100001: out_v[45] = 10'b1000101110;
    16'b0001000000110001: out_v[45] = 10'b1001001011;
    16'b0011000000001001: out_v[45] = 10'b1111100000;
    16'b0000000000100001: out_v[45] = 10'b0001101101;
    16'b0011000000100001: out_v[45] = 10'b0000011110;
    16'b0011000010100001: out_v[45] = 10'b0000011011;
    16'b0011000010110001: out_v[45] = 10'b1110110110;
    16'b0001000010111001: out_v[45] = 10'b0010110001;
    16'b0001000000011001: out_v[45] = 10'b1110010100;
    16'b0001000010110001: out_v[45] = 10'b1011011110;
    16'b0001000000010001: out_v[45] = 10'b0110011011;
    16'b0010000010110001: out_v[45] = 10'b0111011110;
    16'b0000000010100001: out_v[45] = 10'b1001000110;
    16'b0010000010000001: out_v[45] = 10'b1101001000;
    16'b0010000000110001: out_v[45] = 10'b1101100111;
    16'b0001000000000001: out_v[45] = 10'b1001011111;
    16'b0001000010000001: out_v[45] = 10'b0111110101;
    16'b0011000010101001: out_v[45] = 10'b1101001000;
    16'b0011000010100000: out_v[45] = 10'b0001111000;
    16'b0001000000011000: out_v[45] = 10'b1100001000;
    16'b0001000000111011: out_v[45] = 10'b0101111010;
    16'b0001000010110011: out_v[45] = 10'b1111110101;
    16'b0001000000000011: out_v[45] = 10'b0101000110;
    16'b0001000010111011: out_v[45] = 10'b0010110010;
    16'b0001000010101000: out_v[45] = 10'b0111100110;
    16'b0001000010000000: out_v[45] = 10'b0010110110;
    16'b0011000010100010: out_v[45] = 10'b1011100110;
    16'b0001000000101011: out_v[45] = 10'b1001000010;
    16'b0001000010100000: out_v[45] = 10'b0000101001;
    16'b0001000010100010: out_v[45] = 10'b1011100110;
    16'b0001000000110011: out_v[45] = 10'b0001111000;
    16'b0001000010101001: out_v[45] = 10'b0101101000;
    16'b0001000000100011: out_v[45] = 10'b1010100110;
    16'b0001000000011010: out_v[45] = 10'b1001100111;
    16'b0001000000100000: out_v[45] = 10'b1111001011;
    16'b0001000000010011: out_v[45] = 10'b0101010101;
    16'b0001000010010001: out_v[45] = 10'b1111110010;
    16'b0001000010100011: out_v[45] = 10'b0110110111;
    16'b0001000000000000: out_v[45] = 10'b0001101001;
    16'b0001000000110000: out_v[45] = 10'b1000001101;
    16'b0001000000101000: out_v[45] = 10'b0101110101;
    16'b0001000000001000: out_v[45] = 10'b0101011011;
    16'b0010000010101001: out_v[45] = 10'b0101010110;
    16'b0010000000001001: out_v[45] = 10'b1111010110;
    16'b0011000000001000: out_v[45] = 10'b0110100001;
    16'b0010000000001000: out_v[45] = 10'b1011110010;
    16'b0011000000101000: out_v[45] = 10'b1111011000;
    16'b0011000010001001: out_v[45] = 10'b0111110011;
    16'b0010000010001000: out_v[45] = 10'b1111001001;
    16'b0010000010101000: out_v[45] = 10'b1010110011;
    16'b0001000010011001: out_v[45] = 10'b1100100000;
    16'b0011000010011001: out_v[45] = 10'b1100110110;
    16'b0000100010000001: out_v[45] = 10'b0001011001;
    16'b0011000000010001: out_v[45] = 10'b1001101110;
    16'b0011000000100000: out_v[45] = 10'b0011001110;
    16'b0010100010011001: out_v[45] = 10'b0011100101;
    16'b0001000010001001: out_v[45] = 10'b1100100011;
    16'b0011000010010001: out_v[45] = 10'b0110110010;
    16'b0011000000010011: out_v[45] = 10'b1100010111;
    16'b0001000010010000: out_v[45] = 10'b1101000010;
    16'b0001000000010000: out_v[45] = 10'b0110110010;
    16'b0011000010010011: out_v[45] = 10'b0101011001;
    16'b0001000010010011: out_v[45] = 10'b0111111011;
    16'b0011000010110011: out_v[45] = 10'b0010100001;
    16'b0000000010111001: out_v[45] = 10'b0100011011;
    default: out_v[45] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1001000000100101: out_v[46] = 10'b1010110101;
    16'b1000000000100101: out_v[46] = 10'b0101010001;
    16'b0000000000100001: out_v[46] = 10'b1110100101;
    16'b0000000001100001: out_v[46] = 10'b0001111011;
    16'b0000000000100101: out_v[46] = 10'b0100111111;
    16'b0000000000000101: out_v[46] = 10'b0100110011;
    16'b0000000000000001: out_v[46] = 10'b0010000101;
    16'b0000000000000000: out_v[46] = 10'b1000011011;
    16'b0000000101100001: out_v[46] = 10'b1010011011;
    16'b1010000000100101: out_v[46] = 10'b1011011000;
    16'b0001000000100101: out_v[46] = 10'b0010010011;
    16'b0001000000100001: out_v[46] = 10'b0010110110;
    16'b0000000101100000: out_v[46] = 10'b1111100101;
    16'b1000000001100101: out_v[46] = 10'b0011000001;
    16'b0000000000100000: out_v[46] = 10'b0010110110;
    16'b0100000101100000: out_v[46] = 10'b1110110111;
    16'b0101000000100000: out_v[46] = 10'b0100011111;
    16'b1000000101100101: out_v[46] = 10'b0111100101;
    16'b1000000000000101: out_v[46] = 10'b0011100110;
    16'b0101000000100001: out_v[46] = 10'b1110110010;
    16'b1000000000000100: out_v[46] = 10'b1001010111;
    16'b1000000000100100: out_v[46] = 10'b1010001001;
    16'b0000000001100101: out_v[46] = 10'b1110011011;
    16'b0000000101100101: out_v[46] = 10'b1010011011;
    16'b0000000001100000: out_v[46] = 10'b1010011111;
    16'b0001000000100000: out_v[46] = 10'b0110000111;
    16'b1010000000000101: out_v[46] = 10'b1000010000;
    16'b1000000000100001: out_v[46] = 10'b0000101001;
    16'b0010000000000000: out_v[46] = 10'b1101000000;
    16'b0011000000100000: out_v[46] = 10'b0010100010;
    16'b0010000001100000: out_v[46] = 10'b0100110000;
    16'b0010000000100000: out_v[46] = 10'b0100110101;
    16'b0010000100100000: out_v[46] = 10'b0001100010;
    16'b0010000001000000: out_v[46] = 10'b1101101010;
    16'b1010000000000000: out_v[46] = 10'b0111100100;
    16'b1010000000000100: out_v[46] = 10'b0010100110;
    16'b0010000101100000: out_v[46] = 10'b1011111010;
    16'b0110000101100000: out_v[46] = 10'b1111010111;
    16'b1010000101000100: out_v[46] = 10'b0010100101;
    16'b0010000101000000: out_v[46] = 10'b0110110101;
    16'b0010000001000100: out_v[46] = 10'b1110111010;
    16'b0000000001000000: out_v[46] = 10'b1000101010;
    16'b0010000101000100: out_v[46] = 10'b0111011001;
    16'b1100000101100100: out_v[46] = 10'b1010110100;
    16'b1010000101100100: out_v[46] = 10'b0010101100;
    16'b1010000001000100: out_v[46] = 10'b1000000111;
    16'b0110000001000000: out_v[46] = 10'b1011100101;
    16'b1110000000000100: out_v[46] = 10'b0001010100;
    16'b0110000101000100: out_v[46] = 10'b1001001011;
    16'b0010000000000100: out_v[46] = 10'b1110000001;
    16'b1000000101000100: out_v[46] = 10'b1000110100;
    16'b0010000001000001: out_v[46] = 10'b1001000110;
    16'b0110000101000000: out_v[46] = 10'b0101001100;
    16'b1000000001000100: out_v[46] = 10'b1110000001;
    16'b1110000001000100: out_v[46] = 10'b1011100101;
    16'b0110000001100000: out_v[46] = 10'b0010001110;
    16'b0010000000000001: out_v[46] = 10'b0011001001;
    16'b0110000000000000: out_v[46] = 10'b1001111000;
    16'b0000000101000000: out_v[46] = 10'b1100010010;
    16'b1110000101100100: out_v[46] = 10'b0100001011;
    16'b0010000000100001: out_v[46] = 10'b0010011011;
    16'b1110000101000100: out_v[46] = 10'b0010010111;
    16'b0010000000000101: out_v[46] = 10'b1100011100;
    16'b0110000000100000: out_v[46] = 10'b0001110110;
    16'b1001000000100000: out_v[46] = 10'b1010110001;
    16'b1010000101100000: out_v[46] = 10'b1011101010;
    16'b1011000000100100: out_v[46] = 10'b0011010110;
    16'b1000000000100000: out_v[46] = 10'b1111011000;
    16'b1011000000100000: out_v[46] = 10'b1011001101;
    16'b0011000000100001: out_v[46] = 10'b0011001011;
    16'b1001000000100100: out_v[46] = 10'b1001001111;
    16'b1000000101100000: out_v[46] = 10'b0100111000;
    16'b1010000000100100: out_v[46] = 10'b0011011010;
    16'b1001000000100001: out_v[46] = 10'b1001100001;
    16'b1010000001100100: out_v[46] = 10'b1011111010;
    16'b1011000000000000: out_v[46] = 10'b0011100111;
    16'b1111000000100100: out_v[46] = 10'b1100110010;
    16'b0011000000000000: out_v[46] = 10'b1100111101;
    16'b1011000000100101: out_v[46] = 10'b0000010100;
    16'b1011000000000100: out_v[46] = 10'b0101011000;
    16'b1010000000100000: out_v[46] = 10'b0111001111;
    16'b1010000000100001: out_v[46] = 10'b1100000000;
    16'b1000000101100100: out_v[46] = 10'b1000001111;
    16'b1010000001100000: out_v[46] = 10'b0000111011;
    16'b1011000000100001: out_v[46] = 10'b0101110000;
    16'b1010000101100001: out_v[46] = 10'b1000001011;
    16'b1000000101100001: out_v[46] = 10'b1110110100;
    16'b1000000000000000: out_v[46] = 10'b0111110100;
    16'b0010000101100001: out_v[46] = 10'b0110000001;
    16'b1010000101100101: out_v[46] = 10'b1111011100;
    16'b1000000001100000: out_v[46] = 10'b1010100111;
    16'b1000000001100001: out_v[46] = 10'b1100001011;
    16'b0100000101100001: out_v[46] = 10'b0011110010;
    16'b1000000001100100: out_v[46] = 10'b1110110110;
    16'b1010000000000001: out_v[46] = 10'b1000110000;
    16'b0010000000100101: out_v[46] = 10'b1101111000;
    16'b0011000000100101: out_v[46] = 10'b1100100010;
    16'b0011000000100100: out_v[46] = 10'b0101111011;
    16'b0010000000100100: out_v[46] = 10'b0011111000;
    16'b1000000000000001: out_v[46] = 10'b1010101010;
    16'b1011000000000101: out_v[46] = 10'b0101101000;
    16'b1010000001100001: out_v[46] = 10'b1110010011;
    16'b0010000001100001: out_v[46] = 10'b0001011100;
    16'b0001000000000001: out_v[46] = 10'b1101100101;
    16'b1111000000100101: out_v[46] = 10'b1011110011;
    16'b1010000001100101: out_v[46] = 10'b0111000010;
    16'b1010000001000101: out_v[46] = 10'b1011101010;
    16'b0010000101000101: out_v[46] = 10'b1100111011;
    16'b1000000001000101: out_v[46] = 10'b0101001000;
    16'b1010000101000101: out_v[46] = 10'b0110001010;
    16'b0010000001100101: out_v[46] = 10'b1011001110;
    16'b0010000100000000: out_v[46] = 10'b1001110011;
    16'b0010000101000001: out_v[46] = 10'b1011100111;
    16'b0010000001000101: out_v[46] = 10'b0011110011;
    16'b0010000100000101: out_v[46] = 10'b1110100000;
    16'b1010000100000101: out_v[46] = 10'b0111001011;
    16'b0001000010100000: out_v[46] = 10'b0011110001;
    16'b0011000010100000: out_v[46] = 10'b1011100111;
    16'b0000000010000000: out_v[46] = 10'b0011111010;
    16'b0000000010000001: out_v[46] = 10'b0011011110;
    16'b0011000010100001: out_v[46] = 10'b0010111111;
    16'b0010000000000011: out_v[46] = 10'b0001111011;
    16'b0001000010000001: out_v[46] = 10'b1001101111;
    16'b0001000010100001: out_v[46] = 10'b0100011010;
    16'b1011000000000001: out_v[46] = 10'b0111000001;
    16'b0011000000000001: out_v[46] = 10'b1101000011;
    16'b0010000010000101: out_v[46] = 10'b1001100100;
    16'b1011000010100101: out_v[46] = 10'b1111000111;
    16'b1010000010000101: out_v[46] = 10'b1100101011;
    16'b0011000010100101: out_v[46] = 10'b1101010111;
    default: out_v[46] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000010000000010: out_v[47] = 10'b0110010110;
    16'b1000010000000010: out_v[47] = 10'b1010111001;
    16'b0000000000000010: out_v[47] = 10'b0101000111;
    16'b1000000000000010: out_v[47] = 10'b0001100001;
    16'b1000000000000000: out_v[47] = 10'b1110110010;
    16'b0000000000000000: out_v[47] = 10'b0100110110;
    16'b0000000000000011: out_v[47] = 10'b0001110111;
    16'b1000010000000000: out_v[47] = 10'b0010010111;
    16'b0000010000000011: out_v[47] = 10'b1001101110;
    16'b0000010000000000: out_v[47] = 10'b0010011010;
    16'b1000000000000011: out_v[47] = 10'b1000101001;
    16'b0000000000000001: out_v[47] = 10'b0001110010;
    16'b0000001000000010: out_v[47] = 10'b0000001100;
    16'b0000010000000001: out_v[47] = 10'b0100001111;
    16'b0000011000000010: out_v[47] = 10'b0101100110;
    16'b0000000100000001: out_v[47] = 10'b0010011001;
    16'b0000000101000001: out_v[47] = 10'b1011100101;
    16'b0000010100000001: out_v[47] = 10'b1111100000;
    16'b0000000100000000: out_v[47] = 10'b1010010001;
    16'b0000010101000001: out_v[47] = 10'b0100011110;
    16'b0000010100000000: out_v[47] = 10'b0101110010;
    16'b1000000000000001: out_v[47] = 10'b0001110111;
    16'b1000010000000001: out_v[47] = 10'b0101110001;
    16'b0000010001000001: out_v[47] = 10'b1011000111;
    16'b0000000000001010: out_v[47] = 10'b0100100000;
    16'b0000010000001010: out_v[47] = 10'b1111100010;
    16'b0000001000000000: out_v[47] = 10'b1111000101;
    16'b1000000000001010: out_v[47] = 10'b1111100010;
    16'b0000011000000000: out_v[47] = 10'b1000011011;
    16'b0000000000001000: out_v[47] = 10'b0101010111;
    16'b1000010100000000: out_v[47] = 10'b0111001000;
    16'b1000010101000001: out_v[47] = 10'b1101011001;
    16'b0000000001000001: out_v[47] = 10'b1111000101;
    16'b1000010001000000: out_v[47] = 10'b1000100011;
    16'b0000010001000000: out_v[47] = 10'b1111101010;
    16'b1000010001000001: out_v[47] = 10'b1100010111;
    16'b0000000001000000: out_v[47] = 10'b1010011010;
    default: out_v[47] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1100101010100000: out_v[48] = 10'b0001100011;
    16'b1000101010100001: out_v[48] = 10'b1001100101;
    16'b0000100010100000: out_v[48] = 10'b0011100001;
    16'b1100011000100000: out_v[48] = 10'b1111001010;
    16'b1000001000100000: out_v[48] = 10'b0110011111;
    16'b0000000000100000: out_v[48] = 10'b0010110111;
    16'b1000000000101001: out_v[48] = 10'b0110011111;
    16'b1100001000100000: out_v[48] = 10'b1001001101;
    16'b1100111010100000: out_v[48] = 10'b0110110001;
    16'b1100001000101001: out_v[48] = 10'b1001110011;
    16'b1100001000100001: out_v[48] = 10'b0010111101;
    16'b1100110010000000: out_v[48] = 10'b0110000101;
    16'b1000000010101001: out_v[48] = 10'b1101011110;
    16'b1100101010101001: out_v[48] = 10'b0110011111;
    16'b1000001000101000: out_v[48] = 10'b0010111111;
    16'b1100111010100001: out_v[48] = 10'b0110011001;
    16'b1100011010100000: out_v[48] = 10'b1001010110;
    16'b1000101010101001: out_v[48] = 10'b1000011111;
    16'b1100001000000000: out_v[48] = 10'b0111011001;
    16'b1000001000101001: out_v[48] = 10'b1011111110;
    16'b1100101010000000: out_v[48] = 10'b0101110010;
    16'b1000100010101001: out_v[48] = 10'b0000110101;
    16'b1000001010100001: out_v[48] = 10'b0101111011;
    16'b1100010010000000: out_v[48] = 10'b0000001111;
    16'b1100011010000000: out_v[48] = 10'b1100001100;
    16'b0100100010101001: out_v[48] = 10'b0111000011;
    16'b1000101010100000: out_v[48] = 10'b1011000111;
    16'b0000000000101001: out_v[48] = 10'b0001111011;
    16'b0000001000100000: out_v[48] = 10'b0000010111;
    16'b0000101010100000: out_v[48] = 10'b1000110101;
    16'b1000001010101001: out_v[48] = 10'b0101010110;
    16'b1100101000100000: out_v[48] = 10'b1111000110;
    16'b1100101010100001: out_v[48] = 10'b1011100110;
    16'b1000001000100001: out_v[48] = 10'b1110011000;
    16'b1100100010101001: out_v[48] = 10'b1111011011;
    16'b0100110010101001: out_v[48] = 10'b0110010111;
    16'b1100110010101001: out_v[48] = 10'b0111110011;
    16'b1100001010100000: out_v[48] = 10'b0101111110;
    16'b1100011000000000: out_v[48] = 10'b0100110010;
    16'b1100000000000000: out_v[48] = 10'b0110100010;
    16'b1100111010000000: out_v[48] = 10'b0000001011;
    16'b1000101010101000: out_v[48] = 10'b1011011110;
    16'b0100110010000001: out_v[48] = 10'b0010011001;
    16'b0100110010000000: out_v[48] = 10'b0010110111;
    16'b1100001010100001: out_v[48] = 10'b1111010111;
    16'b1000001010100000: out_v[48] = 10'b1111111000;
    16'b0000100010101001: out_v[48] = 10'b0000111001;
    16'b1100001000101000: out_v[48] = 10'b1000110111;
    16'b1000100010000000: out_v[48] = 10'b0111000000;
    16'b0000000000000000: out_v[48] = 10'b0000001011;
    16'b0000000000001000: out_v[48] = 10'b1000001010;
    16'b0000000000000001: out_v[48] = 10'b1010110000;
    16'b0000100000000000: out_v[48] = 10'b1110110101;
    16'b1000100000000000: out_v[48] = 10'b1101011011;
    16'b1000101010000000: out_v[48] = 10'b1101011000;
    16'b0000000000001001: out_v[48] = 10'b1100100101;
    16'b0000101010000000: out_v[48] = 10'b0110000111;
    16'b0000100010000000: out_v[48] = 10'b0101100001;
    16'b1000000000000000: out_v[48] = 10'b0001010011;
    16'b0000100000000001: out_v[48] = 10'b1101000010;
    16'b1000101000001000: out_v[48] = 10'b1110001111;
    16'b1100011010001000: out_v[48] = 10'b1011010110;
    16'b0000100000001000: out_v[48] = 10'b1010010101;
    16'b1000101010001001: out_v[48] = 10'b1010001010;
    16'b1000101010001000: out_v[48] = 10'b0100110010;
    16'b0000100010001001: out_v[48] = 10'b0001111001;
    16'b1000011010001000: out_v[48] = 10'b1000010010;
    16'b0100110010001000: out_v[48] = 10'b1110000110;
    16'b1000110010001000: out_v[48] = 10'b1001110100;
    16'b0000110010001000: out_v[48] = 10'b1110100110;
    16'b1000111010001000: out_v[48] = 10'b1010100010;
    16'b0100111010000000: out_v[48] = 10'b0101011100;
    16'b1000011010000000: out_v[48] = 10'b1001010110;
    16'b0100100010000000: out_v[48] = 10'b0011011110;
    16'b1000001000001000: out_v[48] = 10'b1110011000;
    16'b0000100010001000: out_v[48] = 10'b1011101000;
    16'b1100111010001000: out_v[48] = 10'b0101110100;
    16'b1000011000000000: out_v[48] = 10'b0110110001;
    16'b0000011000001000: out_v[48] = 10'b1111011111;
    16'b0000111010001000: out_v[48] = 10'b1101110001;
    16'b0100100010001000: out_v[48] = 10'b0101101111;
    16'b1100011000001000: out_v[48] = 10'b1110110011;
    16'b1000100010001000: out_v[48] = 10'b0010110101;
    16'b0100111010001000: out_v[48] = 10'b1010110011;
    16'b1000011000001000: out_v[48] = 10'b1101011101;
    16'b0100000000001000: out_v[48] = 10'b0001011101;
    16'b0000101010001000: out_v[48] = 10'b0001110100;
    16'b1000100000001000: out_v[48] = 10'b0101010100;
    16'b0000111010000000: out_v[48] = 10'b0100011110;
    16'b1000111010000000: out_v[48] = 10'b1011011110;
    16'b0100100000001000: out_v[48] = 10'b1100110100;
    16'b1000111010001001: out_v[48] = 10'b0011101011;
    16'b0000011010000000: out_v[48] = 10'b0111011010;
    16'b0100011000000000: out_v[48] = 10'b1111100000;
    16'b0000110010000000: out_v[48] = 10'b1101110010;
    16'b1100110010001000: out_v[48] = 10'b1001000111;
    16'b1000100010001001: out_v[48] = 10'b0111110101;
    16'b0000011000000000: out_v[48] = 10'b0100110111;
    16'b0100011010000000: out_v[48] = 10'b1011101010;
    16'b0100000000000000: out_v[48] = 10'b1101101100;
    16'b1100101010001000: out_v[48] = 10'b1011000001;
    16'b0100010000000000: out_v[48] = 10'b0001001110;
    16'b1100111000001001: out_v[48] = 10'b1101100011;
    16'b0000100010000001: out_v[48] = 10'b0100111100;
    16'b1000111010000001: out_v[48] = 10'b0011101010;
    16'b1100101010001001: out_v[48] = 10'b0011011101;
    16'b0100110000001001: out_v[48] = 10'b1011011011;
    16'b1000011000001001: out_v[48] = 10'b1101110011;
    16'b1000110000001001: out_v[48] = 10'b0101110010;
    16'b1100111010101000: out_v[48] = 10'b0011011110;
    16'b1000010000001001: out_v[48] = 10'b1101001011;
    16'b0100100000001001: out_v[48] = 10'b1000111011;
    16'b1100110000001001: out_v[48] = 10'b1001111010;
    16'b0000100000001001: out_v[48] = 10'b1001101101;
    16'b1100110010001001: out_v[48] = 10'b1111001010;
    16'b1100111010001001: out_v[48] = 10'b0000001111;
    16'b1100100010001001: out_v[48] = 10'b1000111011;
    16'b0100010000001001: out_v[48] = 10'b0000110101;
    16'b1100111010101001: out_v[48] = 10'b1110000011;
    16'b0100000000001001: out_v[48] = 10'b0100011001;
    16'b0100100010000001: out_v[48] = 10'b1111001000;
    16'b0000010000001001: out_v[48] = 10'b0110100000;
    16'b0100100010001001: out_v[48] = 10'b1001101101;
    16'b0100110010001001: out_v[48] = 10'b0110011001;
    16'b1100100010000000: out_v[48] = 10'b0101101000;
    16'b1100111010000001: out_v[48] = 10'b1111011101;
    16'b1000111000001000: out_v[48] = 10'b0011111110;
    16'b1000111000001001: out_v[48] = 10'b1100110111;
    16'b1100010000001001: out_v[48] = 10'b0011111011;
    16'b1100100010001000: out_v[48] = 10'b0011111011;
    16'b1000110010001001: out_v[48] = 10'b1101110101;
    16'b0100110010100001: out_v[48] = 10'b1011110110;
    16'b0100110000100000: out_v[48] = 10'b1100100011;
    16'b0100100000000000: out_v[48] = 10'b0110001101;
    16'b0100010010100000: out_v[48] = 10'b1000110111;
    16'b0100110000100001: out_v[48] = 10'b0101110110;
    16'b0100110010100000: out_v[48] = 10'b0001110010;
    16'b0100110010101000: out_v[48] = 10'b0110011101;
    16'b0100010000100000: out_v[48] = 10'b1100110101;
    16'b1100010000100000: out_v[48] = 10'b1001110111;
    16'b0000110010100000: out_v[48] = 10'b1110110001;
    16'b0100100010100000: out_v[48] = 10'b1001111011;
    16'b0100010010000000: out_v[48] = 10'b0011010011;
    16'b1100010010100000: out_v[48] = 10'b0101110110;
    16'b0100010000101001: out_v[48] = 10'b0010100100;
    16'b0100100010100001: out_v[48] = 10'b0110110001;
    16'b0100100000100000: out_v[48] = 10'b1010000101;
    16'b0100010010100001: out_v[48] = 10'b0000110111;
    16'b0100100000100001: out_v[48] = 10'b1101011100;
    16'b0100010010101001: out_v[48] = 10'b0110110111;
    16'b0000110010100001: out_v[48] = 10'b1011001010;
    16'b0000010010100000: out_v[48] = 10'b1011110010;
    16'b0000010000100000: out_v[48] = 10'b1011101000;
    16'b1100110010100000: out_v[48] = 10'b1010010001;
    16'b0100010000100001: out_v[48] = 10'b1101111100;
    16'b0100010010000001: out_v[48] = 10'b1110011111;
    16'b0100010010101000: out_v[48] = 10'b0011111101;
    16'b0000010010100001: out_v[48] = 10'b0011111010;
    16'b0100100000000001: out_v[48] = 10'b0100111110;
    16'b1100010000101001: out_v[48] = 10'b0111110110;
    16'b1100011000100001: out_v[48] = 10'b1101010010;
    16'b1100001000000001: out_v[48] = 10'b1000010111;
    16'b1100011000101001: out_v[48] = 10'b1110110110;
    16'b0100000000100000: out_v[48] = 10'b0011110101;
    16'b1000001000000000: out_v[48] = 10'b1000110100;
    16'b0000010000101001: out_v[48] = 10'b0100111010;
    16'b1000011000100001: out_v[48] = 10'b1110010110;
    16'b0100000000000001: out_v[48] = 10'b0001110101;
    16'b0100000000101001: out_v[48] = 10'b1010100001;
    16'b1100000000100000: out_v[48] = 10'b0110101110;
    16'b1100100010100000: out_v[48] = 10'b1101111001;
    16'b1100000000100001: out_v[48] = 10'b0100011111;
    16'b0100101010000000: out_v[48] = 10'b1110110010;
    16'b1100000000000001: out_v[48] = 10'b0011001111;
    16'b0100000000100001: out_v[48] = 10'b1011101000;
    16'b1000011000101001: out_v[48] = 10'b1011011111;
    16'b1100000000101001: out_v[48] = 10'b0011111101;
    16'b1100011000001001: out_v[48] = 10'b1000110001;
    16'b1100010000100001: out_v[48] = 10'b0001101101;
    16'b0100101010100000: out_v[48] = 10'b1010111010;
    16'b0100000000000010: out_v[48] = 10'b1001011000;
    16'b0100010000100010: out_v[48] = 10'b0001011111;
    16'b0100010000000010: out_v[48] = 10'b0101001011;
    16'b0100000000101000: out_v[48] = 10'b1110011011;
    16'b0100010000101000: out_v[48] = 10'b1011001000;
    16'b1100010000000000: out_v[48] = 10'b1101011011;
    16'b0000000000000010: out_v[48] = 10'b0011110001;
    16'b0000010000100010: out_v[48] = 10'b1111001001;
    16'b0100010000001000: out_v[48] = 10'b1011001000;
    16'b0000100010101000: out_v[48] = 10'b1011011011;
    16'b0100000000100010: out_v[48] = 10'b0011011100;
    16'b0000010000101000: out_v[48] = 10'b0011011010;
    16'b0100011000100010: out_v[48] = 10'b1101011110;
    16'b0000010000000000: out_v[48] = 10'b1001001111;
    16'b0100011000000010: out_v[48] = 10'b1111001011;
    16'b0100100010101000: out_v[48] = 10'b0101110000;
    16'b1100010000000010: out_v[48] = 10'b0011001000;
    16'b0000000000101000: out_v[48] = 10'b0101011111;
    16'b1100011000100010: out_v[48] = 10'b1011011000;
    16'b1000110010100100: out_v[48] = 10'b0100011100;
    16'b0000100010100001: out_v[48] = 10'b1000101110;
    16'b0000110010100100: out_v[48] = 10'b1001111011;
    16'b0000110010000001: out_v[48] = 10'b0111110010;
    16'b0000100010000100: out_v[48] = 10'b1101100101;
    16'b1000110010000100: out_v[48] = 10'b1101011110;
    16'b0000100010100100: out_v[48] = 10'b0111110001;
    16'b0000110010000100: out_v[48] = 10'b1100110000;
    16'b0100110010100100: out_v[48] = 10'b0001001110;
    16'b0000010010000100: out_v[48] = 10'b0000101111;
    16'b1000110010100000: out_v[48] = 10'b0011001101;
    16'b0000010010000000: out_v[48] = 10'b0010110010;
    16'b1000110010000000: out_v[48] = 10'b1111101010;
    16'b0000010010100100: out_v[48] = 10'b0110110011;
    16'b1000010010000000: out_v[48] = 10'b1010101000;
    16'b1000010000000000: out_v[48] = 10'b0111100110;
    16'b1000101010000001: out_v[48] = 10'b1010011100;
    16'b1100101010000001: out_v[48] = 10'b0011001101;
    16'b1100100010000001: out_v[48] = 10'b1010011111;
    16'b1000000010000000: out_v[48] = 10'b0111010011;
    16'b1100001010000000: out_v[48] = 10'b1111011010;
    16'b1000001010000000: out_v[48] = 10'b0110000001;
    16'b1000100010000001: out_v[48] = 10'b0011010101;
    16'b1100110010100001: out_v[48] = 10'b1011101100;
    16'b1100100010100001: out_v[48] = 10'b0110100110;
    16'b0000110010001001: out_v[48] = 10'b0111001100;
    16'b0100010000100100: out_v[48] = 10'b1001010101;
    16'b0100010010100100: out_v[48] = 10'b1101110111;
    16'b0100100010000100: out_v[48] = 10'b0011101011;
    16'b0100110010000100: out_v[48] = 10'b0110100001;
    16'b0000010000100001: out_v[48] = 10'b1100100110;
    default: out_v[48] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0111001000000000: out_v[49] = 10'b1001110111;
    16'b0011001000000000: out_v[49] = 10'b0100110011;
    16'b0001001000100000: out_v[49] = 10'b0000111101;
    16'b0011001000100000: out_v[49] = 10'b1100000011;
    16'b0001001000000000: out_v[49] = 10'b0011001010;
    16'b0001000000100000: out_v[49] = 10'b0000000011;
    16'b0111000000000000: out_v[49] = 10'b1001100011;
    16'b0000001000000000: out_v[49] = 10'b0111001011;
    16'b0010001000100000: out_v[49] = 10'b1110011000;
    16'b0010000000000000: out_v[49] = 10'b0000011101;
    16'b0101000000000000: out_v[49] = 10'b0010100001;
    16'b0001000000000000: out_v[49] = 10'b0010000111;
    16'b0111001000100000: out_v[49] = 10'b0110110100;
    16'b0101001000100000: out_v[49] = 10'b0011101111;
    16'b0100000000000000: out_v[49] = 10'b0100001001;
    16'b0111000000100000: out_v[49] = 10'b1111010001;
    16'b0010001000000000: out_v[49] = 10'b1100110010;
    16'b0011101000100000: out_v[49] = 10'b0000011001;
    16'b0100000000100000: out_v[49] = 10'b1011001111;
    16'b0011000000000000: out_v[49] = 10'b1100110110;
    16'b0010000000100000: out_v[49] = 10'b1110011100;
    16'b0011001000000100: out_v[49] = 10'b0111100011;
    16'b0101001000000000: out_v[49] = 10'b1010111011;
    16'b0000000000100000: out_v[49] = 10'b0001011111;
    16'b0101000000100000: out_v[49] = 10'b0010110010;
    16'b0110000000100000: out_v[49] = 10'b0010011011;
    16'b0110000000000000: out_v[49] = 10'b0001111011;
    16'b0011000000100000: out_v[49] = 10'b0110100011;
    16'b0000001000100000: out_v[49] = 10'b0000111100;
    16'b0010000000000100: out_v[49] = 10'b0101011110;
    16'b0000000000000100: out_v[49] = 10'b0010110000;
    16'b0000001000000100: out_v[49] = 10'b1101110100;
    16'b0000000000000000: out_v[49] = 10'b1110100100;
    16'b0100001000000100: out_v[49] = 10'b0001001010;
    16'b0000100000000100: out_v[49] = 10'b1101011110;
    16'b0010001000000100: out_v[49] = 10'b0101001011;
    16'b0110001000000100: out_v[49] = 10'b0011100101;
    16'b0100000000000100: out_v[49] = 10'b1001001011;
    16'b0110001000000000: out_v[49] = 10'b0110110110;
    16'b0010000000100100: out_v[49] = 10'b1101100000;
    16'b0110000000000100: out_v[49] = 10'b0100000101;
    16'b0010001000100100: out_v[49] = 10'b1000000100;
    16'b0110001000100100: out_v[49] = 10'b0011001001;
    16'b0110000000100100: out_v[49] = 10'b0001010101;
    16'b0101001000000100: out_v[49] = 10'b1111000110;
    16'b0000000000100100: out_v[49] = 10'b0110100101;
    16'b0011000000100100: out_v[49] = 10'b0111011110;
    16'b0000001000100100: out_v[49] = 10'b0101011010;
    16'b0100001000000000: out_v[49] = 10'b0011111101;
    16'b0001001000000100: out_v[49] = 10'b1101101000;
    16'b0111001000000100: out_v[49] = 10'b0110110111;
    16'b0001000000000100: out_v[49] = 10'b1010011111;
    16'b0011000000000100: out_v[49] = 10'b1010010000;
    16'b0101000000000100: out_v[49] = 10'b0110110000;
    16'b0110001000100000: out_v[49] = 10'b1110110110;
    16'b0001100000000100: out_v[49] = 10'b0000011100;
    16'b0111000000000100: out_v[49] = 10'b0101011011;
    16'b0001101000000100: out_v[49] = 10'b0110100111;
    16'b0111100000000000: out_v[49] = 10'b1101101111;
    16'b0001101000000000: out_v[49] = 10'b1100111110;
    16'b0010101000000100: out_v[49] = 10'b1011100010;
    16'b0011101000000100: out_v[49] = 10'b0110010001;
    16'b0011101000000000: out_v[49] = 10'b0011011111;
    16'b0010101000000000: out_v[49] = 10'b1010101111;
    16'b0001101000100000: out_v[49] = 10'b1101111001;
    16'b0111101000000100: out_v[49] = 10'b0001001011;
    16'b0010101000100000: out_v[49] = 10'b1000110010;
    16'b0000101000000100: out_v[49] = 10'b1110100111;
    16'b0000101000000000: out_v[49] = 10'b1010110100;
    16'b0011001000100100: out_v[49] = 10'b0111000100;
    16'b0001001000100100: out_v[49] = 10'b1001000001;
    16'b0010100000000100: out_v[49] = 10'b1111001010;
    default: out_v[49] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000010000100: out_v[50] = 10'b0000111010;
    16'b1001000000000100: out_v[50] = 10'b1001100011;
    16'b1001000011000100: out_v[50] = 10'b0010111010;
    16'b1000010011000000: out_v[50] = 10'b1001000011;
    16'b1000010011000100: out_v[50] = 10'b0001100111;
    16'b1000000000000100: out_v[50] = 10'b1110110001;
    16'b1000000011000100: out_v[50] = 10'b0000100010;
    16'b1001000001000100: out_v[50] = 10'b0010000111;
    16'b0000000001000100: out_v[50] = 10'b0110100011;
    16'b1000010001000100: out_v[50] = 10'b0100111010;
    16'b1000010010000100: out_v[50] = 10'b1111011101;
    16'b1000010000000100: out_v[50] = 10'b1111100001;
    16'b1000000001000100: out_v[50] = 10'b1110100000;
    16'b1001010000000100: out_v[50] = 10'b1011010110;
    16'b1000000010000000: out_v[50] = 10'b0101001100;
    16'b1000000011000000: out_v[50] = 10'b0111000111;
    16'b1000000010000100: out_v[50] = 10'b0000010011;
    16'b1000010001000000: out_v[50] = 10'b0011001011;
    16'b1000000001000000: out_v[50] = 10'b1111000011;
    16'b1000000011010000: out_v[50] = 10'b1001100100;
    16'b0000000011000100: out_v[50] = 10'b0010001100;
    16'b1000000011010100: out_v[50] = 10'b0011011110;
    16'b1001000011000000: out_v[50] = 10'b0110110011;
    16'b1000010011010000: out_v[50] = 10'b0000110011;
    16'b1001010011000100: out_v[50] = 10'b1011011111;
    16'b0000000011000000: out_v[50] = 10'b1101110101;
    16'b0000000000000100: out_v[50] = 10'b0100110111;
    16'b0000010011000000: out_v[50] = 10'b1101010011;
    16'b1001010001000100: out_v[50] = 10'b0001011001;
    16'b0001000000000100: out_v[50] = 10'b0100110100;
    16'b0100000000000000: out_v[50] = 10'b0011000010;
    16'b1100000000000000: out_v[50] = 10'b0001001110;
    16'b1100010010000000: out_v[50] = 10'b0001101011;
    16'b1100010000000000: out_v[50] = 10'b1000101001;
    16'b1100000000000100: out_v[50] = 10'b1100110000;
    16'b1100000010000000: out_v[50] = 10'b0010011100;
    16'b1100000010000100: out_v[50] = 10'b1101110010;
    16'b0100010000000000: out_v[50] = 10'b1000100111;
    16'b0000000000000000: out_v[50] = 10'b1110101011;
    16'b1100010000000100: out_v[50] = 10'b0111001010;
    16'b1000000000000000: out_v[50] = 10'b1101011001;
    16'b0000010000000000: out_v[50] = 10'b0010111110;
    16'b0101000000000000: out_v[50] = 10'b1011010011;
    16'b0100000010000100: out_v[50] = 10'b0110010010;
    16'b1100010010000100: out_v[50] = 10'b1100100001;
    16'b1100100010010000: out_v[50] = 10'b1011110110;
    16'b1100010010010000: out_v[50] = 10'b1010111011;
    16'b0100000000000100: out_v[50] = 10'b1001011100;
    16'b1000010010000000: out_v[50] = 10'b1010101100;
    16'b1100010000010000: out_v[50] = 10'b1101101111;
    16'b1000010000000000: out_v[50] = 10'b1101000100;
    16'b1100110010010000: out_v[50] = 10'b0111001011;
    16'b0100010010000000: out_v[50] = 10'b1101101000;
    16'b0100010000010000: out_v[50] = 10'b1010110001;
    16'b0000010100000000: out_v[50] = 10'b1110100000;
    16'b0100110000010000: out_v[50] = 10'b1101111101;
    16'b0000010000010000: out_v[50] = 10'b0110011011;
    16'b0100000000010000: out_v[50] = 10'b0100000111;
    16'b0100010100000000: out_v[50] = 10'b0001100111;
    16'b1100000010010000: out_v[50] = 10'b1011101101;
    16'b0000000000010000: out_v[50] = 10'b0001110111;
    16'b0100000001000100: out_v[50] = 10'b0100101100;
    16'b1100000000010000: out_v[50] = 10'b1110101001;
    16'b0100000010000000: out_v[50] = 10'b1000001000;
    16'b0100100000010000: out_v[50] = 10'b0111010110;
    16'b1000010000010000: out_v[50] = 10'b1011110010;
    16'b1000000000010000: out_v[50] = 10'b0011110110;
    16'b0100010000000100: out_v[50] = 10'b0011001010;
    16'b1100100000010000: out_v[50] = 10'b0100100101;
    16'b0000000010000000: out_v[50] = 10'b0010011001;
    16'b1100010110000000: out_v[50] = 10'b1110010111;
    16'b1101000000000000: out_v[50] = 10'b1110101000;
    16'b1100000110000000: out_v[50] = 10'b1000010001;
    16'b1100000011000100: out_v[50] = 10'b0010011000;
    16'b0100000011000000: out_v[50] = 10'b0100010001;
    16'b1100000011000000: out_v[50] = 10'b1101100100;
    16'b1100000100000000: out_v[50] = 10'b1010011111;
    16'b1100010011000100: out_v[50] = 10'b0101001011;
    16'b0100000011000100: out_v[50] = 10'b1000101011;
    16'b1100010100000000: out_v[50] = 10'b1110100011;
    16'b1100000001000100: out_v[50] = 10'b0011001111;
    16'b1101000001000100: out_v[50] = 10'b1100010110;
    16'b1100000001000000: out_v[50] = 10'b1001010001;
    16'b1101000011000000: out_v[50] = 10'b0101110000;
    16'b0101000001000000: out_v[50] = 10'b0001111111;
    16'b1101000001000000: out_v[50] = 10'b1100101110;
    16'b1101000000000100: out_v[50] = 10'b0111000110;
    16'b0100000001000000: out_v[50] = 10'b1101010000;
    16'b0100000001000010: out_v[50] = 10'b0010011010;
    16'b0101000000000100: out_v[50] = 10'b1110011000;
    16'b0101000001000100: out_v[50] = 10'b1000010100;
    16'b0100010011000000: out_v[50] = 10'b0110100011;
    16'b0000000001000000: out_v[50] = 10'b0001110001;
    16'b0001000011000000: out_v[50] = 10'b0101010111;
    16'b1001000001000000: out_v[50] = 10'b0111100000;
    16'b1101000011000100: out_v[50] = 10'b0000010100;
    16'b1001000010000100: out_v[50] = 10'b1000110010;
    16'b0001000011000100: out_v[50] = 10'b1000101101;
    16'b1101000010000100: out_v[50] = 10'b1110100111;
    16'b1100010011000000: out_v[50] = 10'b0111010011;
    16'b0101000011000000: out_v[50] = 10'b0110001001;
    16'b0101000011000100: out_v[50] = 10'b1100000110;
    16'b1100000001010000: out_v[50] = 10'b0111001011;
    16'b1100010001000100: out_v[50] = 10'b0010101111;
    16'b0000010000000100: out_v[50] = 10'b1101000010;
    16'b1100010001000000: out_v[50] = 10'b0000111110;
    16'b1100011000000100: out_v[50] = 10'b0110110111;
    16'b1100001000000100: out_v[50] = 10'b0110110101;
    16'b1000000001001100: out_v[50] = 10'b1001110011;
    16'b0100000000001100: out_v[50] = 10'b1111000101;
    16'b1100000000001100: out_v[50] = 10'b1100101111;
    16'b1100000001001100: out_v[50] = 10'b1100100010;
    16'b1000000000001000: out_v[50] = 10'b0110100101;
    16'b1000000000001100: out_v[50] = 10'b1111000100;
    16'b0100000000001000: out_v[50] = 10'b0110010011;
    16'b1100000001001000: out_v[50] = 10'b1101110101;
    16'b1100000000001000: out_v[50] = 10'b1011000110;
    16'b0100000001001100: out_v[50] = 10'b0011000101;
    16'b1001000001001100: out_v[50] = 10'b1011101111;
    16'b1000000001001000: out_v[50] = 10'b1000010111;
    16'b1101010000000100: out_v[50] = 10'b1111110010;
    16'b0100010010000100: out_v[50] = 10'b0101010001;
    default: out_v[50] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001100000100010: out_v[51] = 10'b1100010001;
    16'b0001000001101010: out_v[51] = 10'b1101110100;
    16'b0000100001101010: out_v[51] = 10'b1001011110;
    16'b0000000001001010: out_v[51] = 10'b0001011001;
    16'b0001000000000010: out_v[51] = 10'b0001011011;
    16'b0001000001100000: out_v[51] = 10'b0000011101;
    16'b0000000001000010: out_v[51] = 10'b0000011110;
    16'b0000000001101000: out_v[51] = 10'b0001101011;
    16'b0000000000100000: out_v[51] = 10'b0010100110;
    16'b0000100001000010: out_v[51] = 10'b1000000111;
    16'b0001000001100010: out_v[51] = 10'b1000110011;
    16'b0000000001101010: out_v[51] = 10'b0011001011;
    16'b0001100001101010: out_v[51] = 10'b0010101011;
    16'b0001000001001010: out_v[51] = 10'b1111000011;
    16'b0001100001000010: out_v[51] = 10'b1000101011;
    16'b0001000000100000: out_v[51] = 10'b1000110111;
    16'b0000000001100010: out_v[51] = 10'b1111011001;
    16'b0001000000100010: out_v[51] = 10'b0001110001;
    16'b0001000001101000: out_v[51] = 10'b0010000110;
    16'b0001100000000010: out_v[51] = 10'b0100101011;
    16'b0000100001001010: out_v[51] = 10'b1000001010;
    16'b0001100001001010: out_v[51] = 10'b1101010101;
    16'b0000100000000010: out_v[51] = 10'b0100011011;
    16'b0000000000000010: out_v[51] = 10'b1010101110;
    16'b0001100001100010: out_v[51] = 10'b1111110000;
    16'b0001000001000010: out_v[51] = 10'b0111100100;
    16'b0100100001001010: out_v[51] = 10'b0000001011;
    16'b0000000001000000: out_v[51] = 10'b1101110001;
    16'b0000000000000000: out_v[51] = 10'b1011100010;
    16'b0010000001000000: out_v[51] = 10'b0010000111;
    16'b0001000001000000: out_v[51] = 10'b0101011011;
    16'b0000100000100010: out_v[51] = 10'b0110100010;
    16'b0001000000000000: out_v[51] = 10'b1010010100;
    16'b0000000001001000: out_v[51] = 10'b1001101101;
    16'b0001000001001000: out_v[51] = 10'b0110100110;
    16'b0000000000100010: out_v[51] = 10'b0111110100;
    16'b0100100000000010: out_v[51] = 10'b0000100101;
    16'b1001000001101000: out_v[51] = 10'b1101100010;
    16'b0000000001100000: out_v[51] = 10'b0100001110;
    16'b1000000001101000: out_v[51] = 10'b1011011111;
    16'b1000000001001010: out_v[51] = 10'b1011100010;
    16'b1001000001100000: out_v[51] = 10'b0010000111;
    16'b1001100001101010: out_v[51] = 10'b1000011100;
    16'b0101100001101010: out_v[51] = 10'b1011010011;
    16'b1001000001001000: out_v[51] = 10'b0011110111;
    16'b0100100001000010: out_v[51] = 10'b0011011101;
    16'b0000000000101000: out_v[51] = 10'b1011000011;
    16'b0001000000001000: out_v[51] = 10'b1111001001;
    16'b1000000001101010: out_v[51] = 10'b0111011011;
    16'b1001000001101010: out_v[51] = 10'b1010111100;
    16'b1001000000100000: out_v[51] = 10'b1001100100;
    16'b1000100001000010: out_v[51] = 10'b1100110011;
    16'b0001000000101000: out_v[51] = 10'b1011000101;
    16'b1001000001100010: out_v[51] = 10'b1110111111;
    16'b0101100001001010: out_v[51] = 10'b1010100110;
    16'b0000100001100010: out_v[51] = 10'b1011111011;
    16'b1000100001001010: out_v[51] = 10'b1101100101;
    16'b1000000001100000: out_v[51] = 10'b1001100001;
    16'b1000000001000010: out_v[51] = 10'b0010010111;
    16'b1001100001001010: out_v[51] = 10'b1110011101;
    16'b0101100000000010: out_v[51] = 10'b0111111010;
    16'b0011000000100010: out_v[51] = 10'b0111111111;
    16'b0010000000100010: out_v[51] = 10'b0000011110;
    16'b0011000000100000: out_v[51] = 10'b1000111111;
    16'b0101100000100010: out_v[51] = 10'b1001011000;
    16'b0101100000000000: out_v[51] = 10'b1101100011;
    16'b0101100000100000: out_v[51] = 10'b1100101011;
    16'b0101000000000000: out_v[51] = 10'b1100100011;
    16'b0100100000100010: out_v[51] = 10'b0010110110;
    16'b0100100000000000: out_v[51] = 10'b1000110101;
    16'b1000000000000010: out_v[51] = 10'b0010110101;
    16'b1001000000100010: out_v[51] = 10'b1101001101;
    16'b1001000000000010: out_v[51] = 10'b1001000001;
    16'b1000000000100000: out_v[51] = 10'b0010011010;
    16'b1001100000100010: out_v[51] = 10'b0011011001;
    16'b1000000000100010: out_v[51] = 10'b1111101101;
    16'b1001100000000010: out_v[51] = 10'b1111000010;
    16'b1001000000000000: out_v[51] = 10'b1000011101;
    16'b0000000000110010: out_v[51] = 10'b1100011111;
    16'b0010010001000000: out_v[51] = 10'b1011000000;
    16'b0010000000000000: out_v[51] = 10'b1101011000;
    16'b0000000000010000: out_v[51] = 10'b1111100101;
    16'b0000000000110000: out_v[51] = 10'b0011000110;
    16'b0000100000100000: out_v[51] = 10'b1101011000;
    16'b0010000001001000: out_v[51] = 10'b1011111010;
    16'b0011000001001000: out_v[51] = 10'b0011110011;
    16'b0001100000000000: out_v[51] = 10'b1101001011;
    16'b0011000001000000: out_v[51] = 10'b1001011000;
    16'b0100000000000000: out_v[51] = 10'b1100111010;
    default: out_v[51] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000011100000: out_v[52] = 10'b0011010001;
    16'b1000000001100000: out_v[52] = 10'b0011010011;
    16'b0100100010100000: out_v[52] = 10'b1111000001;
    16'b0000100011100000: out_v[52] = 10'b1110000110;
    16'b0010000001100000: out_v[52] = 10'b0001111010;
    16'b1010000001100000: out_v[52] = 10'b1101100001;
    16'b0010000001000000: out_v[52] = 10'b1110011000;
    16'b0000000011000000: out_v[52] = 10'b1110110011;
    16'b0110000001000000: out_v[52] = 10'b0000010101;
    16'b1100100011100000: out_v[52] = 10'b0000011111;
    16'b1000000011100000: out_v[52] = 10'b0100110010;
    16'b0000000001100000: out_v[52] = 10'b1000110100;
    16'b0000100010100000: out_v[52] = 10'b1111101011;
    16'b0100100011100000: out_v[52] = 10'b1100110010;
    16'b0110100011100000: out_v[52] = 10'b1101000110;
    16'b0010000011100000: out_v[52] = 10'b0101011011;
    16'b0110100010100000: out_v[52] = 10'b1101101000;
    16'b0100100010000000: out_v[52] = 10'b1010100011;
    16'b1000001001100000: out_v[52] = 10'b1110110101;
    16'b1000000001000000: out_v[52] = 10'b0110001111;
    16'b1100100010000000: out_v[52] = 10'b0110110111;
    16'b1010001001100000: out_v[52] = 10'b1011100111;
    16'b1010000001000000: out_v[52] = 10'b1011001010;
    16'b0010100011100000: out_v[52] = 10'b0011001011;
    16'b0110100010000000: out_v[52] = 10'b0111000100;
    16'b0000000001000000: out_v[52] = 10'b1000110000;
    16'b1100100011000000: out_v[52] = 10'b0011111010;
    16'b0000000010000000: out_v[52] = 10'b1101001110;
    16'b1110100011100000: out_v[52] = 10'b0011001011;
    16'b0110000011100000: out_v[52] = 10'b1101011111;
    16'b0000000010100000: out_v[52] = 10'b0101010111;
    16'b0100100000000000: out_v[52] = 10'b0101111111;
    16'b1010000011100000: out_v[52] = 10'b0110110001;
    16'b0110000001100000: out_v[52] = 10'b0110001111;
    16'b0010000011000000: out_v[52] = 10'b1011110010;
    16'b1000000011000000: out_v[52] = 10'b0101000001;
    16'b1100100010100000: out_v[52] = 10'b0111010010;
    16'b0100100000100000: out_v[52] = 10'b0000010111;
    16'b1010000000000000: out_v[52] = 10'b0001011101;
    16'b0010000000000000: out_v[52] = 10'b0000110111;
    16'b0000000000000000: out_v[52] = 10'b0001011110;
    16'b0010000010000000: out_v[52] = 10'b0110110101;
    16'b1000000000000000: out_v[52] = 10'b1100100010;
    16'b0010100010000000: out_v[52] = 10'b0010110101;
    16'b0010000010100000: out_v[52] = 10'b1011001110;
    16'b0010000000100000: out_v[52] = 10'b0111110100;
    16'b0010100000000000: out_v[52] = 10'b1011010100;
    16'b0010110010000000: out_v[52] = 10'b0001010101;
    16'b1010001010100000: out_v[52] = 10'b0001010111;
    16'b1010000010100000: out_v[52] = 10'b0110011111;
    16'b0010110010100000: out_v[52] = 10'b1000010110;
    16'b0000100000100000: out_v[52] = 10'b0111110011;
    16'b0010100000100000: out_v[52] = 10'b0001011011;
    16'b0010100010100000: out_v[52] = 10'b1011001111;
    16'b0010110000000000: out_v[52] = 10'b1010011001;
    16'b1010100010100000: out_v[52] = 10'b1101110111;
    16'b1010100010000000: out_v[52] = 10'b1011001110;
    16'b0000100010000000: out_v[52] = 10'b1001001010;
    16'b0000000000100000: out_v[52] = 10'b0100110110;
    16'b0000100000000000: out_v[52] = 10'b0111110000;
    16'b1010000000100000: out_v[52] = 10'b0110001101;
    16'b1010101010100000: out_v[52] = 10'b0001101000;
    16'b1010000010000000: out_v[52] = 10'b0110001011;
    16'b1010001000100000: out_v[52] = 10'b0111100100;
    16'b1010001010000000: out_v[52] = 10'b1011111110;
    16'b0010100011000000: out_v[52] = 10'b1100101101;
    16'b1000001000000000: out_v[52] = 10'b1011011011;
    16'b0000110010000000: out_v[52] = 10'b0000101011;
    16'b0000110011000000: out_v[52] = 10'b0001001100;
    16'b0000100011000000: out_v[52] = 10'b1000111001;
    16'b0000110010100000: out_v[52] = 10'b1011101000;
    16'b1000001010000000: out_v[52] = 10'b1001000111;
    16'b0000001010000000: out_v[52] = 10'b1011100101;
    16'b0000110011100000: out_v[52] = 10'b1001001110;
    16'b0000101010000000: out_v[52] = 10'b0011110011;
    16'b1000000010000000: out_v[52] = 10'b1011000001;
    16'b1000101010000000: out_v[52] = 10'b1010010101;
    16'b0000110000000000: out_v[52] = 10'b1010010101;
    16'b1000100010000000: out_v[52] = 10'b1001111111;
    16'b0000100001000000: out_v[52] = 10'b0111110010;
    16'b1000100010100000: out_v[52] = 10'b1000011011;
    16'b0000100001100000: out_v[52] = 10'b0110011000;
    16'b0100000000000000: out_v[52] = 10'b1001111000;
    16'b0100010000000000: out_v[52] = 10'b0001111010;
    16'b1100100000000000: out_v[52] = 10'b0001110101;
    16'b1100100000100000: out_v[52] = 10'b1110011011;
    16'b0100010000100000: out_v[52] = 10'b0110011011;
    16'b1000100000000000: out_v[52] = 10'b0001001010;
    16'b1000100000100000: out_v[52] = 10'b1010101000;
    16'b0100110000100000: out_v[52] = 10'b0010111111;
    16'b0100000000100000: out_v[52] = 10'b1111011000;
    16'b1010000011000000: out_v[52] = 10'b1000111010;
    16'b1110100000100000: out_v[52] = 10'b0110010010;
    16'b1000100011000000: out_v[52] = 10'b1111100001;
    16'b1000100001000000: out_v[52] = 10'b1000100110;
    16'b1000100011100000: out_v[52] = 10'b0011111111;
    16'b1100100001000000: out_v[52] = 10'b1100100011;
    16'b1100000000000000: out_v[52] = 10'b0001111111;
    16'b0110110000100000: out_v[52] = 10'b1001100001;
    16'b0110100000100000: out_v[52] = 10'b0001001000;
    16'b0110100000000000: out_v[52] = 10'b0011010011;
    16'b0010100001100000: out_v[52] = 10'b0111000001;
    16'b0100000001100000: out_v[52] = 10'b1111001000;
    16'b0100000001000000: out_v[52] = 10'b1011001101;
    16'b0010100001000000: out_v[52] = 10'b0100111001;
    16'b0100100001100000: out_v[52] = 10'b0110011110;
    16'b0100110001100000: out_v[52] = 10'b1111010110;
    16'b0000110000100000: out_v[52] = 10'b0111110101;
    16'b0110100001100000: out_v[52] = 10'b0010101001;
    16'b0110000000000000: out_v[52] = 10'b1101101111;
    16'b0010110000100000: out_v[52] = 10'b0110000101;
    16'b0100100001000000: out_v[52] = 10'b1100110101;
    16'b1110100010000000: out_v[52] = 10'b0110010011;
    16'b1010100011000000: out_v[52] = 10'b1101001001;
    16'b1010100011100000: out_v[52] = 10'b0001000110;
    16'b0100100010100010: out_v[52] = 10'b1101000111;
    16'b0110000000100000: out_v[52] = 10'b1000111010;
    16'b0100000010000000: out_v[52] = 10'b0011111010;
    16'b0100100010000010: out_v[52] = 10'b1010001101;
    16'b0100000010100000: out_v[52] = 10'b0101101010;
    default: out_v[52] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000001000001100: out_v[53] = 10'b0011010001;
    16'b1000000000011111: out_v[53] = 10'b1011011111;
    16'b1000000000011010: out_v[53] = 10'b1001001111;
    16'b1000000000010110: out_v[53] = 10'b0010001001;
    16'b1000001000001100: out_v[53] = 10'b1111011000;
    16'b1000000000010100: out_v[53] = 10'b1000100011;
    16'b1000000000011000: out_v[53] = 10'b0001110011;
    16'b0000000000010110: out_v[53] = 10'b0111011011;
    16'b1000000000010000: out_v[53] = 10'b0000110001;
    16'b1000000000011100: out_v[53] = 10'b1101011010;
    16'b1000001000011110: out_v[53] = 10'b0101000000;
    16'b1000000000011110: out_v[53] = 10'b0011001001;
    16'b1000001000001110: out_v[53] = 10'b1100000011;
    16'b0000000000011110: out_v[53] = 10'b0100011101;
    16'b1000001000011100: out_v[53] = 10'b0010110010;
    16'b1000001000011010: out_v[53] = 10'b0111001011;
    16'b1000000000001110: out_v[53] = 10'b1100001110;
    16'b0000000000000100: out_v[53] = 10'b1011000101;
    16'b0000000000011111: out_v[53] = 10'b1010110110;
    16'b1000000000000100: out_v[53] = 10'b1011111011;
    16'b0000000000001010: out_v[53] = 10'b0111110011;
    16'b1000000000000000: out_v[53] = 10'b0011100100;
    16'b0000000000001000: out_v[53] = 10'b0100010110;
    16'b1000001000011111: out_v[53] = 10'b0100000011;
    16'b0000000000001110: out_v[53] = 10'b1011000110;
    16'b0000000000000110: out_v[53] = 10'b1111110101;
    16'b1000000010010100: out_v[53] = 10'b0011110011;
    16'b1000001000011000: out_v[53] = 10'b0011111010;
    16'b1000000000001100: out_v[53] = 10'b1000101100;
    16'b0000000000001100: out_v[53] = 10'b1100100001;
    16'b0000001000000010: out_v[53] = 10'b1000101010;
    16'b0000000000000010: out_v[53] = 10'b1100010011;
    16'b0000000000000000: out_v[53] = 10'b0010011010;
    16'b1000001000000010: out_v[53] = 10'b1111111010;
    16'b0000001000000100: out_v[53] = 10'b1110000010;
    16'b1000000000000010: out_v[53] = 10'b1101111111;
    16'b1000001000010000: out_v[53] = 10'b0000101111;
    16'b1000001000000011: out_v[53] = 10'b1111011111;
    16'b0000000000000011: out_v[53] = 10'b0111010011;
    16'b0000001000000000: out_v[53] = 10'b1001110100;
    16'b1000001000000000: out_v[53] = 10'b0101001101;
    16'b1000001000000100: out_v[53] = 10'b0011101110;
    16'b1000001000010100: out_v[53] = 10'b1001010111;
    16'b1000000000000110: out_v[53] = 10'b0000011100;
    16'b1000001000010110: out_v[53] = 10'b0111010100;
    16'b0000001000010100: out_v[53] = 10'b0101110110;
    16'b0000000010000100: out_v[53] = 10'b0001010111;
    16'b1000011000010100: out_v[53] = 10'b0011100101;
    16'b1000001000000110: out_v[53] = 10'b0111001000;
    16'b1000010000010100: out_v[53] = 10'b1111011010;
    16'b0000001000000111: out_v[53] = 10'b0001011011;
    16'b0000001000001110: out_v[53] = 10'b0000111010;
    16'b0000001000001111: out_v[53] = 10'b1000011010;
    16'b0000000010001110: out_v[53] = 10'b1101100011;
    16'b0000001000000110: out_v[53] = 10'b1010111010;
    16'b0000001010001100: out_v[53] = 10'b0100011011;
    16'b0000001010001110: out_v[53] = 10'b1100010001;
    16'b0000001010001111: out_v[53] = 10'b1011111000;
    16'b0000000000000111: out_v[53] = 10'b0000010001;
    16'b0000001010000100: out_v[53] = 10'b0110111000;
    16'b0000000000001111: out_v[53] = 10'b1011110000;
    16'b0000000010001100: out_v[53] = 10'b1101110011;
    16'b0000001000001000: out_v[53] = 10'b1000110101;
    16'b0000001000001011: out_v[53] = 10'b1001101100;
    16'b0000011000000000: out_v[53] = 10'b0010110001;
    16'b0000001000001010: out_v[53] = 10'b1000110000;
    16'b0000011010000000: out_v[53] = 10'b0110111001;
    16'b0000001010001000: out_v[53] = 10'b0110001111;
    16'b1000001000001000: out_v[53] = 10'b0100011001;
    16'b0000001010000000: out_v[53] = 10'b0011110000;
    16'b1000000000001000: out_v[53] = 10'b1100100111;
    16'b0000000000001011: out_v[53] = 10'b0011100000;
    16'b0000000100001000: out_v[53] = 10'b0100011110;
    16'b0000000010000000: out_v[53] = 10'b1001011010;
    16'b0000000100000000: out_v[53] = 10'b1000001101;
    16'b0000000110001000: out_v[53] = 10'b1011011011;
    16'b0000000110000000: out_v[53] = 10'b0100010110;
    16'b0000000010000011: out_v[53] = 10'b0011110011;
    16'b0000000010001000: out_v[53] = 10'b1000001011;
    16'b0000000010000010: out_v[53] = 10'b0011100111;
    16'b1000001000010111: out_v[53] = 10'b1111000110;
    16'b1000001000001111: out_v[53] = 10'b0101110001;
    16'b1000000000001111: out_v[53] = 10'b0110010111;
    16'b1000001000001010: out_v[53] = 10'b1011100010;
    16'b1000001000011011: out_v[53] = 10'b0001000011;
    16'b0000011000000100: out_v[53] = 10'b1110101010;
    default: out_v[53] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001000000000010: out_v[54] = 10'b0100001000;
    16'b0001000000000011: out_v[54] = 10'b0100001111;
    16'b1001000000000011: out_v[54] = 10'b1101010111;
    16'b0000000000000000: out_v[54] = 10'b0010111010;
    16'b0000000000000010: out_v[54] = 10'b0110010110;
    16'b0000000000000011: out_v[54] = 10'b0010111110;
    16'b1000010000000001: out_v[54] = 10'b1011001111;
    16'b0000010000000011: out_v[54] = 10'b0001111001;
    16'b0001000000000001: out_v[54] = 10'b1000100001;
    16'b0000000000000001: out_v[54] = 10'b0011110001;
    16'b1000000000000001: out_v[54] = 10'b0001010111;
    16'b0001010000000010: out_v[54] = 10'b0011010010;
    16'b0001010000000001: out_v[54] = 10'b1101011011;
    16'b0001000000000000: out_v[54] = 10'b1000100001;
    16'b1000000000000011: out_v[54] = 10'b1110010110;
    16'b0000010000000010: out_v[54] = 10'b0000001111;
    16'b0001010000000011: out_v[54] = 10'b0011111011;
    16'b1001000000000001: out_v[54] = 10'b0100000011;
    16'b0000010000000001: out_v[54] = 10'b0101100000;
    16'b1001010000000001: out_v[54] = 10'b1101010100;
    16'b1000010000000011: out_v[54] = 10'b0110011101;
    16'b0001010000000000: out_v[54] = 10'b0000011110;
    16'b1001010000000011: out_v[54] = 10'b0111110011;
    16'b0000010000000000: out_v[54] = 10'b0101001010;
    16'b0000010000001000: out_v[54] = 10'b1100000101;
    16'b0000000000001010: out_v[54] = 10'b1101011100;
    16'b0001010000001010: out_v[54] = 10'b1100000101;
    16'b1000010000000000: out_v[54] = 10'b0000110110;
    16'b1000010000000010: out_v[54] = 10'b0101001110;
    16'b0000010000001010: out_v[54] = 10'b0111010111;
    16'b0001000000001010: out_v[54] = 10'b0000001100;
    16'b1000000000000010: out_v[54] = 10'b1010101011;
    16'b1001000000000010: out_v[54] = 10'b1000101000;
    16'b0000000000001000: out_v[54] = 10'b1000111010;
    16'b1001000000000000: out_v[54] = 10'b0100100001;
    16'b1001010000000010: out_v[54] = 10'b0011100011;
    16'b1000000000000000: out_v[54] = 10'b0100101001;
    16'b0000000000001011: out_v[54] = 10'b0010011000;
    16'b0000000000001001: out_v[54] = 10'b0001111011;
    16'b0001000000001000: out_v[54] = 10'b1001100111;
    16'b0000010000010000: out_v[54] = 10'b0111000000;
    16'b0000010000010010: out_v[54] = 10'b1111100001;
    16'b0000010000010011: out_v[54] = 10'b1111011001;
    16'b0000010000010001: out_v[54] = 10'b1011001111;
    16'b0000000000000110: out_v[54] = 10'b0010011000;
    default: out_v[54] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000100001010000: out_v[55] = 10'b1010101011;
    16'b0010100001011010: out_v[55] = 10'b1011110110;
    16'b0010100101011010: out_v[55] = 10'b1001001101;
    16'b0010100001010000: out_v[55] = 10'b1001100010;
    16'b0010100001010010: out_v[55] = 10'b1010110001;
    16'b0010100001001000: out_v[55] = 10'b0101100010;
    16'b0011100001011010: out_v[55] = 10'b0000101011;
    16'b0010100101000000: out_v[55] = 10'b1101001111;
    16'b0010000001000000: out_v[55] = 10'b0010111000;
    16'b0010100001000010: out_v[55] = 10'b0011011011;
    16'b0010100001011000: out_v[55] = 10'b0110101011;
    16'b0010100000010000: out_v[55] = 10'b0101100001;
    16'b0000000001010000: out_v[55] = 10'b0010100101;
    16'b0010000001010000: out_v[55] = 10'b1001001001;
    16'b0000100001010010: out_v[55] = 10'b0111100110;
    16'b0110100001010000: out_v[55] = 10'b1110110101;
    16'b0010100001000000: out_v[55] = 10'b0101000010;
    16'b0010000001001000: out_v[55] = 10'b0111100100;
    16'b0011100001010010: out_v[55] = 10'b1000110110;
    16'b0000000001000000: out_v[55] = 10'b1100011111;
    16'b0000100001011000: out_v[55] = 10'b1111000011;
    16'b0010000001011010: out_v[55] = 10'b1010011011;
    16'b0001100001010000: out_v[55] = 10'b1000011111;
    16'b0010100101011000: out_v[55] = 10'b1101011110;
    16'b0011100000011010: out_v[55] = 10'b0011011101;
    16'b0010000001011000: out_v[55] = 10'b1001001011;
    16'b0010000101000000: out_v[55] = 10'b0111000110;
    16'b0010100101010010: out_v[55] = 10'b1111101111;
    16'b0010100101010000: out_v[55] = 10'b1111111101;
    16'b0010100001001010: out_v[55] = 10'b1100100010;
    16'b0010000001010010: out_v[55] = 10'b0011100110;
    16'b0010100101001000: out_v[55] = 10'b0101011011;
    16'b0010000001001010: out_v[55] = 10'b1111110001;
    16'b0000100001000000: out_v[55] = 10'b0001111111;
    16'b0011000001001000: out_v[55] = 10'b0110110010;
    16'b0001000001001000: out_v[55] = 10'b0010010111;
    16'b0000000000001000: out_v[55] = 10'b0111011001;
    16'b0001000000001000: out_v[55] = 10'b1000111100;
    16'b0011000000001000: out_v[55] = 10'b1011010011;
    16'b0000000000001010: out_v[55] = 10'b0001010101;
    16'b0000100000000010: out_v[55] = 10'b0011110011;
    16'b0000000001001000: out_v[55] = 10'b0001001111;
    16'b0000000000000010: out_v[55] = 10'b1111000111;
    16'b0001100000001010: out_v[55] = 10'b1000100011;
    16'b0000100000001010: out_v[55] = 10'b0111011100;
    16'b0001000001001010: out_v[55] = 10'b0011000101;
    16'b0011000000000000: out_v[55] = 10'b1010100010;
    16'b0001000000001010: out_v[55] = 10'b0011111001;
    16'b0000000000000000: out_v[55] = 10'b0101001110;
    16'b0001000000000000: out_v[55] = 10'b0100001111;
    16'b0000000001001010: out_v[55] = 10'b0001001101;
    16'b0001100001001010: out_v[55] = 10'b0110010110;
    16'b0011000001001010: out_v[55] = 10'b0101001001;
    16'b0110000001010010: out_v[55] = 10'b1010000101;
    16'b0011000001000000: out_v[55] = 10'b1100110100;
    16'b0111000000000010: out_v[55] = 10'b1001101000;
    16'b0010000001000010: out_v[55] = 10'b0011011010;
    16'b0111000001001000: out_v[55] = 10'b1110001101;
    16'b0111000001010010: out_v[55] = 10'b0100110111;
    16'b0001000001000010: out_v[55] = 10'b0100000000;
    16'b0111000001000010: out_v[55] = 10'b0010111101;
    16'b0011000000000010: out_v[55] = 10'b0000000101;
    16'b0011000001000010: out_v[55] = 10'b0110011010;
    16'b0011000000010010: out_v[55] = 10'b0100010110;
    16'b0111000000010010: out_v[55] = 10'b1110100100;
    16'b0001000000000010: out_v[55] = 10'b0011101110;
    16'b0011000000010000: out_v[55] = 10'b0010111101;
    16'b0111000000001010: out_v[55] = 10'b1010111111;
    16'b0111000001001010: out_v[55] = 10'b0100010110;
    16'b0011100000001010: out_v[55] = 10'b1011100110;
    16'b0011000000001010: out_v[55] = 10'b1011010100;
    16'b0011000001010010: out_v[55] = 10'b0110110110;
    16'b0011100001000010: out_v[55] = 10'b1111000110;
    16'b0001100000000010: out_v[55] = 10'b1000011000;
    16'b0110000001000010: out_v[55] = 10'b1111100110;
    16'b0011000000011010: out_v[55] = 10'b0010011111;
    16'b0111000001000000: out_v[55] = 10'b0001111100;
    16'b0011100000000010: out_v[55] = 10'b0001001111;
    16'b0001000000011010: out_v[55] = 10'b1101001011;
    16'b0111000000000000: out_v[55] = 10'b1000100101;
    16'b0011000001011010: out_v[55] = 10'b0001101011;
    16'b0001000000010000: out_v[55] = 10'b1100100111;
    16'b0011100000010010: out_v[55] = 10'b0000100101;
    16'b0001000001000000: out_v[55] = 10'b1111010001;
    16'b0011100001000000: out_v[55] = 10'b0110100011;
    16'b0011100000000000: out_v[55] = 10'b0101010101;
    16'b0000000001011000: out_v[55] = 10'b1100011001;
    16'b0010000000001000: out_v[55] = 10'b1111111010;
    16'b0000000001011010: out_v[55] = 10'b1100011110;
    16'b0000000001000010: out_v[55] = 10'b1000111101;
    16'b0000100001001010: out_v[55] = 10'b1001101001;
    16'b0010000000011000: out_v[55] = 10'b0110001010;
    16'b0000000000011000: out_v[55] = 10'b1101001001;
    16'b0000100001001000: out_v[55] = 10'b1111101100;
    16'b0110000001011000: out_v[55] = 10'b1111001000;
    16'b0000100001000010: out_v[55] = 10'b1010100011;
    16'b0000000000011010: out_v[55] = 10'b0111000111;
    16'b0001000000010010: out_v[55] = 10'b0001101010;
    16'b0001100001000010: out_v[55] = 10'b0110011011;
    16'b0000000000010010: out_v[55] = 10'b0110110010;
    16'b0000000000010000: out_v[55] = 10'b1000110100;
    16'b0001100001000000: out_v[55] = 10'b0101001011;
    16'b0001100001010010: out_v[55] = 10'b1100101110;
    16'b0000100000011010: out_v[55] = 10'b0110111000;
    16'b0000100000010000: out_v[55] = 10'b0110010011;
    16'b0001100000010010: out_v[55] = 10'b0101111011;
    16'b0000000000110000: out_v[55] = 10'b0011110011;
    16'b0000100000010010: out_v[55] = 10'b0110010101;
    16'b0000000000110010: out_v[55] = 10'b1100111001;
    16'b0000000001010010: out_v[55] = 10'b1100000110;
    16'b0000100000000000: out_v[55] = 10'b1000101001;
    16'b0001100000011010: out_v[55] = 10'b1011111000;
    16'b0001000001010000: out_v[55] = 10'b0010111101;
    16'b0001100001011000: out_v[55] = 10'b0111010011;
    16'b0001100000010000: out_v[55] = 10'b1000101010;
    16'b0001100000000000: out_v[55] = 10'b0101001011;
    16'b0001100001011010: out_v[55] = 10'b1110010011;
    16'b0010100000000010: out_v[55] = 10'b0111001000;
    16'b0011100001001010: out_v[55] = 10'b0100111100;
    16'b0010100000001010: out_v[55] = 10'b0111010111;
    16'b0010000000001010: out_v[55] = 10'b0111100000;
    16'b0011100001001000: out_v[55] = 10'b1010001111;
    16'b0101100000010010: out_v[55] = 10'b1110100001;
    16'b0101000000000000: out_v[55] = 10'b1111100000;
    16'b0101100001010010: out_v[55] = 10'b0110101111;
    16'b0101100001000010: out_v[55] = 10'b1001011110;
    16'b0111100001010010: out_v[55] = 10'b1010111111;
    16'b0100100001010000: out_v[55] = 10'b0000001011;
    16'b0101100000010000: out_v[55] = 10'b1111011111;
    16'b0110100000010010: out_v[55] = 10'b1101101010;
    16'b0101100001010000: out_v[55] = 10'b0001111111;
    16'b0101100001011010: out_v[55] = 10'b1110100000;
    16'b0101100000000010: out_v[55] = 10'b1100101001;
    16'b0101100001000000: out_v[55] = 10'b0011011110;
    16'b0100100000010010: out_v[55] = 10'b1111101000;
    16'b0111100000010010: out_v[55] = 10'b1101110011;
    16'b0101000000010000: out_v[55] = 10'b1101010001;
    16'b0011100001010000: out_v[55] = 10'b0101000011;
    16'b0101100000000000: out_v[55] = 10'b0011101001;
    16'b0101000000010010: out_v[55] = 10'b0111010001;
    16'b0101000000000010: out_v[55] = 10'b0110011000;
    16'b0100100000010000: out_v[55] = 10'b1110100010;
    16'b0000100000111000: out_v[55] = 10'b1100001110;
    16'b0000110000011010: out_v[55] = 10'b0111100011;
    16'b0001100001001000: out_v[55] = 10'b0111000111;
    16'b0000100000011000: out_v[55] = 10'b1111101000;
    16'b0000100001101010: out_v[55] = 10'b0111101010;
    16'b0000100001011010: out_v[55] = 10'b0010001101;
    16'b0011100000001000: out_v[55] = 10'b0011000101;
    16'b0000110000001010: out_v[55] = 10'b1001101101;
    16'b0000100001111010: out_v[55] = 10'b1111010111;
    16'b0001000001011000: out_v[55] = 10'b0110000000;
    16'b0000100000101010: out_v[55] = 10'b0101110111;
    16'b0000100000111010: out_v[55] = 10'b0111100001;
    16'b0000100000001000: out_v[55] = 10'b1001100101;
    default: out_v[55] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001011000000000: out_v[56] = 10'b0100001111;
    16'b0001010100010000: out_v[56] = 10'b1001001110;
    16'b0001010001010000: out_v[56] = 10'b0111000011;
    16'b0000000101010000: out_v[56] = 10'b0100101110;
    16'b0001010101010000: out_v[56] = 10'b1011111000;
    16'b0000000101010100: out_v[56] = 10'b0111000011;
    16'b0000000100010000: out_v[56] = 10'b1110100101;
    16'b0001010000010000: out_v[56] = 10'b1100000111;
    16'b0000000101000000: out_v[56] = 10'b0001111101;
    16'b0101011000010000: out_v[56] = 10'b1010100110;
    16'b0001000101010000: out_v[56] = 10'b1000001111;
    16'b0101010000010000: out_v[56] = 10'b0110100010;
    16'b0001011000010000: out_v[56] = 10'b0110100001;
    16'b0001011001010000: out_v[56] = 10'b0011110111;
    16'b0101011101010000: out_v[56] = 10'b1010011101;
    16'b0001011101010000: out_v[56] = 10'b1000111111;
    16'b0001010101000000: out_v[56] = 10'b0010100001;
    16'b0101011001010000: out_v[56] = 10'b1010111110;
    16'b0101011001000000: out_v[56] = 10'b0001111000;
    16'b0101010101010000: out_v[56] = 10'b0010101101;
    16'b0001000100010000: out_v[56] = 10'b0011011110;
    16'b0101011000000000: out_v[56] = 10'b1001101001;
    16'b0001010101010100: out_v[56] = 10'b1001101001;
    16'b0001010000000000: out_v[56] = 10'b0111001000;
    16'b0000000001010000: out_v[56] = 10'b0100100001;
    16'b0001010100000000: out_v[56] = 10'b1000100001;
    16'b0000000000010000: out_v[56] = 10'b1100101001;
    16'b0001010001000000: out_v[56] = 10'b1001011101;
    16'b0000000001010100: out_v[56] = 10'b0010010111;
    16'b0001000000010000: out_v[56] = 10'b0110010111;
    16'b0101010001010000: out_v[56] = 10'b0110110110;
    16'b0000000001000100: out_v[56] = 10'b0010100011;
    16'b0001010000000100: out_v[56] = 10'b1111000110;
    16'b0001010001000100: out_v[56] = 10'b1010101010;
    16'b0000000001000000: out_v[56] = 10'b0000011011;
    16'b0000000000000000: out_v[56] = 10'b1011010011;
    16'b0001010100000100: out_v[56] = 10'b1000101000;
    16'b0000000000000100: out_v[56] = 10'b0001011100;
    16'b0001000001000100: out_v[56] = 10'b1000100100;
    16'b0001010101000100: out_v[56] = 10'b0100100110;
    16'b0001000100000100: out_v[56] = 10'b0001111010;
    16'b0001011100000100: out_v[56] = 10'b0110000011;
    16'b0001000000000100: out_v[56] = 10'b0110000000;
    16'b0000000100000100: out_v[56] = 10'b0000111101;
    16'b0101011001000100: out_v[56] = 10'b0101110101;
    16'b0101011101000100: out_v[56] = 10'b0010111111;
    16'b0101010101000100: out_v[56] = 10'b1010011011;
    16'b0101010101000000: out_v[56] = 10'b1100011011;
    16'b0000000000010100: out_v[56] = 10'b1001011101;
    16'b0101010101100100: out_v[56] = 10'b1110100101;
    16'b0001011001000000: out_v[56] = 10'b0010110100;
    16'b0001011101010100: out_v[56] = 10'b0101011010;
    16'b0001010100010100: out_v[56] = 10'b1000111110;
    16'b0100000101000100: out_v[56] = 10'b1001100110;
    16'b0001010000010100: out_v[56] = 10'b1100001010;
    16'b0101011001100100: out_v[56] = 10'b1100010111;
    16'b0101010001000100: out_v[56] = 10'b0110110100;
    16'b0101010100000100: out_v[56] = 10'b1000101000;
    16'b0001011101000100: out_v[56] = 10'b0101110110;
    16'b0100000001000100: out_v[56] = 10'b1011100001;
    16'b0101010001000101: out_v[56] = 10'b0111001001;
    16'b0001011001000100: out_v[56] = 10'b0001010100;
    16'b0101010101010100: out_v[56] = 10'b1000010110;
    16'b0101010101000101: out_v[56] = 10'b0100001001;
    16'b0101000101000100: out_v[56] = 10'b1010100011;
    16'b0101011101100100: out_v[56] = 10'b1001111110;
    16'b0000000101000100: out_v[56] = 10'b1111011100;
    16'b0101011101000000: out_v[56] = 10'b0001010110;
    16'b0001000101000100: out_v[56] = 10'b1101001011;
    16'b0101010101000001: out_v[56] = 10'b0010110011;
    16'b0001010001010100: out_v[56] = 10'b1101110000;
    16'b0101010001010100: out_v[56] = 10'b0110000101;
    16'b0101011000000100: out_v[56] = 10'b1111001100;
    16'b0101010000000100: out_v[56] = 10'b1011000001;
    16'b0101000000000000: out_v[56] = 10'b1100001001;
    16'b0101010100000000: out_v[56] = 10'b0110110110;
    16'b0101010000000000: out_v[56] = 10'b0101011010;
    16'b0101011000100000: out_v[56] = 10'b0110000111;
    16'b0101011000110000: out_v[56] = 10'b1010100001;
    16'b0101010100010000: out_v[56] = 10'b1010100111;
    16'b0101011001100000: out_v[56] = 10'b1001101010;
    16'b0000000100000000: out_v[56] = 10'b0010001001;
    16'b0100000000000000: out_v[56] = 10'b1101110111;
    16'b0101010001000000: out_v[56] = 10'b1100010011;
    16'b0001000101000000: out_v[56] = 10'b0011011011;
    16'b0001000100000000: out_v[56] = 10'b0011011001;
    16'b1101011000100000: out_v[56] = 10'b1101011010;
    16'b0101011100000100: out_v[56] = 10'b0011001011;
    16'b0101001000000000: out_v[56] = 10'b0111011001;
    16'b0101011000100100: out_v[56] = 10'b1001001011;
    16'b0000001100010100: out_v[56] = 10'b0101111111;
    16'b0100001100010000: out_v[56] = 10'b0110001101;
    16'b0000001000010000: out_v[56] = 10'b1010101010;
    16'b0100001000010100: out_v[56] = 10'b0000011010;
    16'b0100000100010100: out_v[56] = 10'b0011111110;
    16'b0100000001010100: out_v[56] = 10'b1001001110;
    16'b0000000100010100: out_v[56] = 10'b1000110110;
    16'b0100000100010000: out_v[56] = 10'b0111010111;
    16'b0000001100010000: out_v[56] = 10'b0011001001;
    16'b0000001000010100: out_v[56] = 10'b1001100010;
    16'b0100000000010000: out_v[56] = 10'b0010011111;
    16'b0001000100010100: out_v[56] = 10'b0000110110;
    16'b0100000000010100: out_v[56] = 10'b0000011111;
    16'b0001000001010100: out_v[56] = 10'b1111000110;
    16'b0100001100010100: out_v[56] = 10'b1010111010;
    16'b0100001000010000: out_v[56] = 10'b0001111100;
    16'b0001011100010100: out_v[56] = 10'b0011100110;
    16'b0001001000010000: out_v[56] = 10'b0001011101;
    16'b0001011000010100: out_v[56] = 10'b1100100000;
    16'b0100000101010100: out_v[56] = 10'b1001100000;
    16'b0001000001000000: out_v[56] = 10'b1110110011;
    16'b0100000101010000: out_v[56] = 10'b0011110010;
    16'b0100000001010000: out_v[56] = 10'b1001001110;
    16'b0001011001010100: out_v[56] = 10'b0111000010;
    16'b0001000101010100: out_v[56] = 10'b1011010111;
    16'b0000001000000000: out_v[56] = 10'b1011101010;
    16'b0000001000100000: out_v[56] = 10'b0001011101;
    16'b1000000100100100: out_v[56] = 10'b0111011011;
    16'b0000000100100000: out_v[56] = 10'b1101101000;
    16'b0000000100100100: out_v[56] = 10'b1111100011;
    16'b1000000100100000: out_v[56] = 10'b1000000100;
    16'b0000001100000000: out_v[56] = 10'b1111110100;
    16'b0100000100000000: out_v[56] = 10'b0011010101;
    16'b0000000001100100: out_v[56] = 10'b1011000000;
    16'b1000001000100000: out_v[56] = 10'b0110010100;
    16'b0000000101100100: out_v[56] = 10'b0101111110;
    16'b0000000000100100: out_v[56] = 10'b0011001101;
    16'b0010000001000100: out_v[56] = 10'b1001010100;
    16'b1000001100100000: out_v[56] = 10'b1111100001;
    16'b0101011001010100: out_v[56] = 10'b0100101010;
    16'b0001011000000100: out_v[56] = 10'b1101011001;
    16'b0101011000010100: out_v[56] = 10'b0110001001;
    16'b0101011101010100: out_v[56] = 10'b0011001111;
    16'b0001011100010000: out_v[56] = 10'b1111000101;
    16'b0101011100010100: out_v[56] = 10'b1101111001;
    default: out_v[56] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0011001000100000: out_v[57] = 10'b1010011011;
    16'b0010001000100010: out_v[57] = 10'b0010011001;
    16'b0010001000000010: out_v[57] = 10'b0110001000;
    16'b0011000000000000: out_v[57] = 10'b0111000101;
    16'b0011000000100000: out_v[57] = 10'b0011010111;
    16'b0010000000100000: out_v[57] = 10'b1001010001;
    16'b0011000000000010: out_v[57] = 10'b1100100101;
    16'b0001000000100000: out_v[57] = 10'b1000111100;
    16'b0110001000100010: out_v[57] = 10'b1011000011;
    16'b0011000000100010: out_v[57] = 10'b0110100101;
    16'b0110001000000010: out_v[57] = 10'b1001101111;
    16'b0001000000000000: out_v[57] = 10'b1011011011;
    16'b0011001000000000: out_v[57] = 10'b0011010111;
    16'b0000001000000010: out_v[57] = 10'b0111011110;
    16'b0011000010100000: out_v[57] = 10'b0010000101;
    16'b0011000010000000: out_v[57] = 10'b0111010111;
    16'b0001001000000010: out_v[57] = 10'b1001101000;
    16'b0001001000100010: out_v[57] = 10'b1010110111;
    16'b0010001000100000: out_v[57] = 10'b0011110010;
    16'b0010000000000000: out_v[57] = 10'b1110110010;
    16'b0001000000000010: out_v[57] = 10'b0111100001;
    16'b0111001000100010: out_v[57] = 10'b0110110000;
    16'b0011001000100010: out_v[57] = 10'b0001000111;
    16'b0010000010100000: out_v[57] = 10'b1000000101;
    16'b0011001000000010: out_v[57] = 10'b0001100100;
    16'b0000001000100010: out_v[57] = 10'b1101111011;
    16'b0001000000100010: out_v[57] = 10'b0110111010;
    16'b0111001000000010: out_v[57] = 10'b1101011011;
    16'b0000000000000000: out_v[57] = 10'b0011010011;
    16'b0100001000100010: out_v[57] = 10'b1001100011;
    16'b0000000000100000: out_v[57] = 10'b1100110101;
    16'b0001001000100000: out_v[57] = 10'b0000110001;
    16'b0011000010100010: out_v[57] = 10'b1100010111;
    16'b0010000000000010: out_v[57] = 10'b0000010100;
    16'b0000001000100000: out_v[57] = 10'b1001011011;
    16'b0110000000000010: out_v[57] = 10'b1100011010;
    16'b0100000000000010: out_v[57] = 10'b0000110011;
    16'b0101001000000010: out_v[57] = 10'b1101001011;
    16'b0100001000000010: out_v[57] = 10'b1110101100;
    16'b0100000000100010: out_v[57] = 10'b0000100110;
    16'b0101000000000010: out_v[57] = 10'b1001011001;
    16'b0101001000000000: out_v[57] = 10'b0111100011;
    16'b0100000000100000: out_v[57] = 10'b1110101110;
    16'b0110000000100010: out_v[57] = 10'b1100110100;
    16'b0100000000000000: out_v[57] = 10'b1001001110;
    16'b0100001000000000: out_v[57] = 10'b0110001011;
    16'b0111000010000010: out_v[57] = 10'b0000100011;
    16'b0111000000100000: out_v[57] = 10'b0011001110;
    16'b0111000000000010: out_v[57] = 10'b1110010001;
    16'b0110000000100000: out_v[57] = 10'b0110100100;
    16'b0010000010000000: out_v[57] = 10'b0010011011;
    16'b0000000010100000: out_v[57] = 10'b0010110000;
    16'b0111000010100010: out_v[57] = 10'b0010011010;
    16'b0001000010100000: out_v[57] = 10'b0110001011;
    16'b0101000000100010: out_v[57] = 10'b1010010101;
    16'b0111000000000000: out_v[57] = 10'b1000101000;
    16'b0101000000100000: out_v[57] = 10'b0100101100;
    16'b0101001000100010: out_v[57] = 10'b0100010000;
    16'b0111000000100010: out_v[57] = 10'b1011110110;
    16'b0110000000000000: out_v[57] = 10'b1100101001;
    16'b0101000000000000: out_v[57] = 10'b0001011010;
    16'b0111001010100010: out_v[57] = 10'b1010001101;
    16'b0000000000100010: out_v[57] = 10'b0100011100;
    16'b0110000010100010: out_v[57] = 10'b0010110111;
    16'b0111000010100000: out_v[57] = 10'b1101101110;
    16'b0011000010000010: out_v[57] = 10'b1101110100;
    16'b0101000010100010: out_v[57] = 10'b0110100110;
    16'b0110000010000010: out_v[57] = 10'b0011010100;
    16'b0101001010100010: out_v[57] = 10'b1101100000;
    16'b0111000010000000: out_v[57] = 10'b0011110010;
    16'b0101001010000010: out_v[57] = 10'b0010001101;
    16'b0101000010000010: out_v[57] = 10'b1100100111;
    16'b0001001010000010: out_v[57] = 10'b1000100010;
    16'b0111001010000010: out_v[57] = 10'b0010001000;
    16'b0110001000000000: out_v[57] = 10'b1001110100;
    16'b0100000010000010: out_v[57] = 10'b0100011011;
    16'b0101000010100000: out_v[57] = 10'b1001101011;
    16'b0101000010000000: out_v[57] = 10'b0001101000;
    16'b0111001000000000: out_v[57] = 10'b0100100100;
    16'b0110001010000010: out_v[57] = 10'b1111100001;
    16'b0100001010000010: out_v[57] = 10'b1011110111;
    16'b0100000010000000: out_v[57] = 10'b1101110010;
    16'b0000000000000010: out_v[57] = 10'b0011111111;
    16'b0010001000000000: out_v[57] = 10'b0011011110;
    16'b0000000010000000: out_v[57] = 10'b1101000111;
    16'b0100000010100000: out_v[57] = 10'b0011010111;
    16'b0001001000000000: out_v[57] = 10'b0000010011;
    16'b0111001010000000: out_v[57] = 10'b0110100010;
    16'b0111001000100000: out_v[57] = 10'b1100110010;
    16'b0110001000100000: out_v[57] = 10'b0110110010;
    16'b0100001000100000: out_v[57] = 10'b1111101101;
    16'b0000001000000000: out_v[57] = 10'b1101010001;
    16'b0000001001000010: out_v[57] = 10'b0111001011;
    16'b0001000001000000: out_v[57] = 10'b0111110101;
    16'b0001000011000010: out_v[57] = 10'b1101110001;
    16'b0000001010000010: out_v[57] = 10'b1111101011;
    16'b0001000010000010: out_v[57] = 10'b0101101101;
    16'b0001000001000010: out_v[57] = 10'b0110111110;
    16'b0000000001000010: out_v[57] = 10'b1110111110;
    16'b0010000010000010: out_v[57] = 10'b1001111100;
    16'b0000000011000010: out_v[57] = 10'b1100010011;
    16'b0000000010000010: out_v[57] = 10'b1111000001;
    16'b0000000001000000: out_v[57] = 10'b0111111101;
    16'b0001000010000000: out_v[57] = 10'b0111101001;
    16'b0001000011000000: out_v[57] = 10'b1100110101;
    16'b0101001000100000: out_v[57] = 10'b0101010001;
    16'b0101000001000000: out_v[57] = 10'b1101100010;
    16'b0100000001000000: out_v[57] = 10'b1101000111;
    16'b0001000000101000: out_v[57] = 10'b1001100111;
    16'b0101000001000010: out_v[57] = 10'b1101110111;
    16'b0100000001000010: out_v[57] = 10'b1001101101;
    16'b0001000001100000: out_v[57] = 10'b1011100011;
    default: out_v[57] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000110001000: out_v[58] = 10'b0100110101;
    16'b1000000010000000: out_v[58] = 10'b1100100011;
    16'b1000000110000000: out_v[58] = 10'b0101110101;
    16'b0000000110000000: out_v[58] = 10'b1001001011;
    16'b0000000000010000: out_v[58] = 10'b1110000101;
    16'b0000000010010000: out_v[58] = 10'b1000110010;
    16'b0000000000000000: out_v[58] = 10'b0011000001;
    16'b0000000010000000: out_v[58] = 10'b0101110001;
    16'b1000000011000000: out_v[58] = 10'b0000010111;
    16'b0000000110010000: out_v[58] = 10'b1111110001;
    16'b0000100110010000: out_v[58] = 10'b0111110101;
    16'b0000000010001000: out_v[58] = 10'b0010110110;
    16'b1000000011010000: out_v[58] = 10'b0001001001;
    16'b1000000110010000: out_v[58] = 10'b1010011101;
    16'b1010000011000000: out_v[58] = 10'b0001100100;
    16'b1000000010010000: out_v[58] = 10'b1010011100;
    16'b1000000000000000: out_v[58] = 10'b0010101011;
    16'b0000000110011000: out_v[58] = 10'b0000001111;
    16'b1010000011001000: out_v[58] = 10'b1010111010;
    16'b0000000100010000: out_v[58] = 10'b1111000001;
    16'b1010000010001000: out_v[58] = 10'b0101011001;
    16'b1000000111000000: out_v[58] = 10'b0000110111;
    16'b1000000010001000: out_v[58] = 10'b1101100111;
    16'b0000000011000000: out_v[58] = 10'b0010110011;
    16'b1000000111010000: out_v[58] = 10'b0000111100;
    16'b0000000010011000: out_v[58] = 10'b0001011111;
    16'b1000000110001000: out_v[58] = 10'b1011000111;
    16'b0000100000010000: out_v[58] = 10'b0000101111;
    16'b0000100010011000: out_v[58] = 10'b1101010010;
    16'b1000100000000000: out_v[58] = 10'b0111001010;
    16'b0000100000000000: out_v[58] = 10'b1101011101;
    16'b0000100010010000: out_v[58] = 10'b0000011111;
    16'b1010100000010000: out_v[58] = 10'b0101001100;
    16'b0010100010010000: out_v[58] = 10'b0111011101;
    16'b0010100000000000: out_v[58] = 10'b0101011010;
    16'b0000100100010000: out_v[58] = 10'b1110100111;
    16'b0000100010000000: out_v[58] = 10'b1001100000;
    16'b0000100000011000: out_v[58] = 10'b0011011111;
    16'b1010100000000000: out_v[58] = 10'b0011111011;
    16'b1000100010010000: out_v[58] = 10'b1010011101;
    16'b1000100000010000: out_v[58] = 10'b1100000110;
    16'b1000100011010000: out_v[58] = 10'b0000011011;
    16'b1000100111000000: out_v[58] = 10'b0110100110;
    16'b0000100001010000: out_v[58] = 10'b0001001110;
    16'b1000100110010000: out_v[58] = 10'b0111000110;
    16'b1000100110000000: out_v[58] = 10'b1110000100;
    16'b1000100100000000: out_v[58] = 10'b0001011000;
    16'b0000100100000000: out_v[58] = 10'b0100011101;
    16'b1000100111010000: out_v[58] = 10'b0100011010;
    16'b1000100010000000: out_v[58] = 10'b1110000000;
    16'b1000100011010100: out_v[58] = 10'b1110000011;
    16'b0000100110000000: out_v[58] = 10'b1111000110;
    16'b1000100011000000: out_v[58] = 10'b0011100011;
    16'b1000100001000000: out_v[58] = 10'b0011101100;
    16'b1000100111010100: out_v[58] = 10'b1011110111;
    16'b1000100001010000: out_v[58] = 10'b1101100111;
    16'b1000100101010000: out_v[58] = 10'b1101011100;
    16'b1000100101000000: out_v[58] = 10'b1111001110;
    16'b1000100100010000: out_v[58] = 10'b0110110100;
    16'b1010000011011000: out_v[58] = 10'b1111011100;
    16'b1000100111011000: out_v[58] = 10'b1101100111;
    16'b1010100011010000: out_v[58] = 10'b0010100011;
    16'b1010000111011000: out_v[58] = 10'b1110010101;
    16'b1010000011010000: out_v[58] = 10'b1011101110;
    16'b0000100110011000: out_v[58] = 10'b1100001110;
    16'b1000000010011000: out_v[58] = 10'b1001011101;
    16'b1000000011011000: out_v[58] = 10'b1101001010;
    16'b1010100111011000: out_v[58] = 10'b1111110111;
    16'b1010100111010000: out_v[58] = 10'b0001001110;
    16'b1010100011011000: out_v[58] = 10'b1010001111;
    16'b1000100011011000: out_v[58] = 10'b0010110011;
    16'b0000100111011000: out_v[58] = 10'b0011101011;
    16'b1000000111011000: out_v[58] = 10'b1101110010;
    16'b1000000001010000: out_v[58] = 10'b1000111100;
    16'b1000100010011000: out_v[58] = 10'b0011001101;
    16'b1000100110011000: out_v[58] = 10'b1011011101;
    16'b0000100110001000: out_v[58] = 10'b1110101010;
    16'b1000000110011000: out_v[58] = 10'b1111011010;
    16'b1000100111001000: out_v[58] = 10'b1101111010;
    16'b1000000001000000: out_v[58] = 10'b1010101101;
    16'b1000000000010000: out_v[58] = 10'b0010101101;
    16'b0010100110010000: out_v[58] = 10'b0001011111;
    16'b0000100100011000: out_v[58] = 10'b1011011110;
    16'b0000100111010001: out_v[58] = 10'b0001011011;
    16'b0010100111010000: out_v[58] = 10'b1110010101;
    16'b0010100100010000: out_v[58] = 10'b1100001001;
    16'b0000100100001000: out_v[58] = 10'b1101010111;
    16'b0000100101010000: out_v[58] = 10'b0001010100;
    16'b0010100101000000: out_v[58] = 10'b0110011010;
    16'b0010100100000000: out_v[58] = 10'b0001010011;
    16'b1010100100010000: out_v[58] = 10'b0001110101;
    16'b1010100101000000: out_v[58] = 10'b1010010101;
    16'b0000100110010001: out_v[58] = 10'b0011011011;
    16'b0010000100000000: out_v[58] = 10'b0111111110;
    16'b0000100101000001: out_v[58] = 10'b0011011110;
    16'b0000100101010001: out_v[58] = 10'b1111101110;
    16'b1010100100000000: out_v[58] = 10'b0010011001;
    16'b0010100101010000: out_v[58] = 10'b0110001101;
    16'b0000100100000001: out_v[58] = 10'b1011010111;
    16'b0000000100000000: out_v[58] = 10'b1000111100;
    16'b1010100110010000: out_v[58] = 10'b0110110100;
    16'b0000100101000000: out_v[58] = 10'b1001011010;
    16'b0000100111010000: out_v[58] = 10'b0110011010;
    16'b1000000100000000: out_v[58] = 10'b1000011110;
    16'b0010100110001000: out_v[58] = 10'b0110101000;
    16'b0000100000110000: out_v[58] = 10'b0011111001;
    16'b1010100111000000: out_v[58] = 10'b0000101100;
    16'b0000100100110000: out_v[58] = 10'b0100001001;
    16'b0000000100110000: out_v[58] = 10'b1010101110;
    16'b0010100110000000: out_v[58] = 10'b1111000111;
    16'b1000100110001000: out_v[58] = 10'b1011101010;
    16'b0000100010001000: out_v[58] = 10'b0011110100;
    16'b1010100111001000: out_v[58] = 10'b1001110011;
    16'b0000000100011000: out_v[58] = 10'b1001100110;
    16'b1010100110001000: out_v[58] = 10'b0100110011;
    16'b0010000110001000: out_v[58] = 10'b1011110001;
    16'b1000100010001000: out_v[58] = 10'b1111001011;
    16'b1000000100010000: out_v[58] = 10'b1101001101;
    16'b1000100101000010: out_v[58] = 10'b0100100111;
    16'b1000100100000010: out_v[58] = 10'b0111101010;
    16'b1000000100000010: out_v[58] = 10'b0100010011;
    16'b1000100000000010: out_v[58] = 10'b1011100011;
    16'b0000100001000000: out_v[58] = 10'b0011011011;
    16'b1000100001000010: out_v[58] = 10'b1111101001;
    16'b1000000101010000: out_v[58] = 10'b1011110000;
    16'b0000100011011000: out_v[58] = 10'b0101011011;
    16'b0010000100010000: out_v[58] = 10'b0010101000;
    16'b0010000000010000: out_v[58] = 10'b0011000010;
    16'b0000100000001000: out_v[58] = 10'b0001011011;
    16'b0010100000010000: out_v[58] = 10'b1011100001;
    16'b0010100011010000: out_v[58] = 10'b1010110001;
    16'b0000000000011000: out_v[58] = 10'b1011100001;
    16'b0010000000010001: out_v[58] = 10'b1100100011;
    16'b0000000000010001: out_v[58] = 10'b1111010000;
    16'b0000100011010000: out_v[58] = 10'b0110110001;
    16'b0000100011001000: out_v[58] = 10'b1110111011;
    16'b0010000000000000: out_v[58] = 10'b0110001011;
    16'b0010100001010000: out_v[58] = 10'b0010101001;
    16'b0000000000001000: out_v[58] = 10'b0111010100;
    16'b0000100001011000: out_v[58] = 10'b1000111011;
    16'b0010100110011000: out_v[58] = 10'b0111010100;
    16'b1010100010000000: out_v[58] = 10'b1011100011;
    16'b1010100110000000: out_v[58] = 10'b1111100110;
    16'b1010100010010000: out_v[58] = 10'b1101000111;
    16'b1000100011001000: out_v[58] = 10'b1111011010;
    16'b1010100011000000: out_v[58] = 10'b1101100011;
    16'b0010100010001000: out_v[58] = 10'b1111100111;
    16'b0010100010000000: out_v[58] = 10'b1111010111;
    16'b0010100110010001: out_v[58] = 10'b1011001001;
    16'b0000100100010001: out_v[58] = 10'b1000100011;
    16'b0010100100010001: out_v[58] = 10'b1100111111;
    default: out_v[58] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000001100000001: out_v[59] = 10'b1101011010;
    16'b0000101100000001: out_v[59] = 10'b0100100000;
    16'b0100001100000001: out_v[59] = 10'b0000110101;
    16'b0000001000000001: out_v[59] = 10'b0100000011;
    16'b0000001100000000: out_v[59] = 10'b0111010100;
    16'b0000101000000001: out_v[59] = 10'b1011000101;
    16'b0000000100000000: out_v[59] = 10'b1010000101;
    16'b0100000000000001: out_v[59] = 10'b1101001010;
    16'b0000000000000001: out_v[59] = 10'b0011010101;
    16'b0000000100000001: out_v[59] = 10'b0010010000;
    16'b0100001000000001: out_v[59] = 10'b0000100110;
    16'b0100000100000001: out_v[59] = 10'b1001001010;
    16'b0100101100000001: out_v[59] = 10'b0001110110;
    16'b0100001000000000: out_v[59] = 10'b0001011101;
    16'b0000001000000000: out_v[59] = 10'b1010101000;
    16'b0100000000000000: out_v[59] = 10'b0110100101;
    16'b0000100100000001: out_v[59] = 10'b0001100010;
    16'b0000100100000000: out_v[59] = 10'b0011100111;
    16'b0000101100000000: out_v[59] = 10'b0000011011;
    16'b0100101000000001: out_v[59] = 10'b0000111011;
    16'b0000000000000000: out_v[59] = 10'b0000111011;
    16'b0100001100000000: out_v[59] = 10'b0100100110;
    16'b0100000100000000: out_v[59] = 10'b0100100010;
    16'b0000001101000001: out_v[59] = 10'b1011011100;
    16'b0000001101000000: out_v[59] = 10'b0001001010;
    16'b0100001101000001: out_v[59] = 10'b0110001110;
    16'b0000100000000000: out_v[59] = 10'b0110101000;
    16'b1000100000000000: out_v[59] = 10'b1011101100;
    16'b0000101000000000: out_v[59] = 10'b0100010110;
    16'b0000100000000001: out_v[59] = 10'b0100011011;
    16'b0001001100000001: out_v[59] = 10'b0010110101;
    16'b0001001100000000: out_v[59] = 10'b1101001011;
    16'b0001001000000001: out_v[59] = 10'b1011100010;
    16'b0001000100000001: out_v[59] = 10'b1111001110;
    16'b0001000100000000: out_v[59] = 10'b1101001011;
    16'b0000000100010001: out_v[59] = 10'b1111000111;
    16'b0000001100010001: out_v[59] = 10'b1100001011;
    16'b0000001000010001: out_v[59] = 10'b1101001010;
    default: out_v[59] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010000000010000: out_v[60] = 10'b0101000001;
    16'b0010101000000010: out_v[60] = 10'b1001101010;
    16'b0000100000110010: out_v[60] = 10'b1000000100;
    16'b0000101010010010: out_v[60] = 10'b0100010011;
    16'b0010001000010000: out_v[60] = 10'b0000000001;
    16'b0000100000000010: out_v[60] = 10'b1111010001;
    16'b0000100000010010: out_v[60] = 10'b1001010011;
    16'b0000101000000010: out_v[60] = 10'b0101010010;
    16'b0010000000000000: out_v[60] = 10'b1101000101;
    16'b0010101010010010: out_v[60] = 10'b0110010100;
    16'b0010100000010010: out_v[60] = 10'b0110110110;
    16'b0000101010000010: out_v[60] = 10'b1101011001;
    16'b0000101000010010: out_v[60] = 10'b1000001001;
    16'b0000000000000000: out_v[60] = 10'b0100010110;
    16'b0000000000010000: out_v[60] = 10'b0010111000;
    16'b0000100000010000: out_v[60] = 10'b0011111100;
    16'b0010100000010000: out_v[60] = 10'b0000111100;
    16'b0000101000110010: out_v[60] = 10'b0101011011;
    16'b0000100000000000: out_v[60] = 10'b1111000010;
    16'b0000001000010000: out_v[60] = 10'b0100001100;
    16'b0010101000010010: out_v[60] = 10'b0111010100;
    16'b0000101000010000: out_v[60] = 10'b1100001111;
    16'b0000101000100010: out_v[60] = 10'b0101110011;
    16'b0010001000000000: out_v[60] = 10'b1001100011;
    16'b0000100000100010: out_v[60] = 10'b1000000011;
    16'b0000100010010010: out_v[60] = 10'b1101010111;
    16'b0010101000010000: out_v[60] = 10'b1010011110;
    16'b0000000000110010: out_v[60] = 10'b1101000001;
    16'b0010101010000010: out_v[60] = 10'b1110001111;
    16'b0000101000000000: out_v[60] = 10'b1001000100;
    16'b0000001000000000: out_v[60] = 10'b0110110000;
    16'b0010001010010000: out_v[60] = 10'b0000011101;
    16'b0010000010010000: out_v[60] = 10'b0111011010;
    16'b0010100000000010: out_v[60] = 10'b0111010100;
    16'b0010001010000000: out_v[60] = 10'b1001110001;
    16'b0010000000000010: out_v[60] = 10'b0110010111;
    16'b0000001010010000: out_v[60] = 10'b1000001100;
    16'b0000000000000010: out_v[60] = 10'b0001101100;
    16'b0001000000000000: out_v[60] = 10'b1000011101;
    16'b0000000000100000: out_v[60] = 10'b0110001100;
    16'b0000001000010010: out_v[60] = 10'b0001011010;
    16'b0010000000010010: out_v[60] = 10'b1111100000;
    16'b0010001000010010: out_v[60] = 10'b0010011111;
    16'b0000000010000000: out_v[60] = 10'b1110010011;
    16'b0011000000000000: out_v[60] = 10'b0010100110;
    16'b0010001000000010: out_v[60] = 10'b1010011100;
    16'b0000001010010010: out_v[60] = 10'b1011001000;
    16'b0000001010000000: out_v[60] = 10'b1101100010;
    16'b0010001010010010: out_v[60] = 10'b1100000111;
    16'b0010000000001000: out_v[60] = 10'b1000000110;
    16'b0010100000000000: out_v[60] = 10'b1101111000;
    16'b0010001010000010: out_v[60] = 10'b1110011011;
    16'b0000000010010000: out_v[60] = 10'b0101110011;
    16'b0010000010000000: out_v[60] = 10'b1101011000;
    16'b0010101010010000: out_v[60] = 10'b1011001110;
    16'b0011100000000000: out_v[60] = 10'b0010101011;
    16'b0001000001000000: out_v[60] = 10'b0110001101;
    16'b0000001000000010: out_v[60] = 10'b0010100000;
    16'b0010101000000000: out_v[60] = 10'b0001101100;
    16'b0010100000110010: out_v[60] = 10'b0001110010;
    16'b0010100000110000: out_v[60] = 10'b1100000011;
    16'b0010100000100000: out_v[60] = 10'b1101010011;
    16'b0000000000010010: out_v[60] = 10'b1001110100;
    16'b0000001000100000: out_v[60] = 10'b1001111110;
    16'b0010001000000100: out_v[60] = 10'b1011111010;
    16'b0000000000110000: out_v[60] = 10'b0011010011;
    16'b0000000100110000: out_v[60] = 10'b0010010001;
    16'b0000000100100000: out_v[60] = 10'b0011010110;
    16'b0000100000110000: out_v[60] = 10'b1110101101;
    16'b0001000000010000: out_v[60] = 10'b0001000100;
    16'b0001000100110000: out_v[60] = 10'b1001101110;
    16'b0000000100000000: out_v[60] = 10'b1001011111;
    16'b0010000000110000: out_v[60] = 10'b0111001010;
    16'b0010100000100010: out_v[60] = 10'b0011111001;
    16'b0000100000100000: out_v[60] = 10'b0111001010;
    default: out_v[60] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1100110100001000: out_v[61] = 10'b0100111111;
    16'b0000000100001000: out_v[61] = 10'b1000010101;
    16'b0001001100001100: out_v[61] = 10'b0000011010;
    16'b1100010100001000: out_v[61] = 10'b1010011011;
    16'b0001101110001101: out_v[61] = 10'b1001011110;
    16'b1100110110001000: out_v[61] = 10'b1010100011;
    16'b0001001101001101: out_v[61] = 10'b0100000011;
    16'b1110110100001000: out_v[61] = 10'b0110111101;
    16'b0010000100001000: out_v[61] = 10'b0001010111;
    16'b0100010100001000: out_v[61] = 10'b0100110011;
    16'b0000100110001000: out_v[61] = 10'b1101010001;
    16'b0001001100001000: out_v[61] = 10'b1001010111;
    16'b0001101110001100: out_v[61] = 10'b0010010111;
    16'b1101110100001000: out_v[61] = 10'b1010010011;
    16'b0100110100001000: out_v[61] = 10'b1001110111;
    16'b0110010000001000: out_v[61] = 10'b0010010111;
    16'b0001100110001100: out_v[61] = 10'b0111011110;
    16'b1110110000001000: out_v[61] = 10'b1100111100;
    16'b0001101111001101: out_v[61] = 10'b1111100001;
    16'b0000100100001000: out_v[61] = 10'b0111111011;
    16'b0000010100001000: out_v[61] = 10'b1100011001;
    16'b0001101011001101: out_v[61] = 10'b1000001011;
    16'b0000001100001000: out_v[61] = 10'b1011001011;
    16'b0000110100001000: out_v[61] = 10'b1111111100;
    16'b0000000100001100: out_v[61] = 10'b0010010111;
    16'b0001001101001100: out_v[61] = 10'b1100000001;
    16'b1000110100001000: out_v[61] = 10'b1111000011;
    16'b1101110100001101: out_v[61] = 10'b1111111110;
    16'b1100110100001101: out_v[61] = 10'b0010011111;
    16'b1100110100001100: out_v[61] = 10'b0100010111;
    16'b0000000011001101: out_v[61] = 10'b1100101101;
    16'b0000000001001001: out_v[61] = 10'b1001010011;
    16'b0011000100000001: out_v[61] = 10'b1001011010;
    16'b0010000000000101: out_v[61] = 10'b0101110011;
    16'b0001000100000101: out_v[61] = 10'b1001000110;
    16'b0001000101000101: out_v[61] = 10'b0010000011;
    16'b0000000000000001: out_v[61] = 10'b0000001001;
    16'b0000000001000101: out_v[61] = 10'b1010100100;
    16'b0000000000000101: out_v[61] = 10'b0011100110;
    16'b0001000100000001: out_v[61] = 10'b0011000001;
    16'b0000000011001001: out_v[61] = 10'b1111001011;
    16'b0011000001000101: out_v[61] = 10'b0111001110;
    16'b0000000001000001: out_v[61] = 10'b1100100111;
    16'b0000000001001101: out_v[61] = 10'b1000101011;
    16'b0001001101000101: out_v[61] = 10'b1111001001;
    16'b0011000101000101: out_v[61] = 10'b0111000100;
    16'b0000000010001000: out_v[61] = 10'b1100001010;
    16'b0011000100000101: out_v[61] = 10'b0101001111;
    16'b0001001001001101: out_v[61] = 10'b1001101101;
    16'b0000000000001001: out_v[61] = 10'b0100110011;
    16'b0001000000000101: out_v[61] = 10'b0000100110;
    16'b0000000011001000: out_v[61] = 10'b1011001011;
    16'b0001000001000101: out_v[61] = 10'b0101110101;
    16'b0000000000001000: out_v[61] = 10'b0011001001;
    16'b0001000000000001: out_v[61] = 10'b1100110111;
    16'b0001000001001101: out_v[61] = 10'b1010011011;
    16'b0001001100000101: out_v[61] = 10'b0110001110;
    16'b0011000000000001: out_v[61] = 10'b1111110101;
    16'b0010000001000101: out_v[61] = 10'b0001011110;
    16'b0011000000000101: out_v[61] = 10'b1100100101;
    16'b0010000000000001: out_v[61] = 10'b1101100111;
    16'b0000000000000000: out_v[61] = 10'b0010100100;
    16'b0000000101000101: out_v[61] = 10'b0010101110;
    16'b0000000001001000: out_v[61] = 10'b1101000110;
    16'b0001001000001000: out_v[61] = 10'b0110100111;
    16'b0001001001001000: out_v[61] = 10'b1010000100;
    16'b0101011101001000: out_v[61] = 10'b1110110101;
    16'b0000000101001001: out_v[61] = 10'b1011110111;
    16'b0001011000001000: out_v[61] = 10'b1001100100;
    16'b0101011001000000: out_v[61] = 10'b0001000111;
    16'b0001001101001000: out_v[61] = 10'b0100011100;
    16'b0101011001001000: out_v[61] = 10'b0000011011;
    16'b0001001000000000: out_v[61] = 10'b1010100000;
    16'b0101011000001000: out_v[61] = 10'b0100101110;
    16'b0101010101001101: out_v[61] = 10'b1010100101;
    16'b0001001001000000: out_v[61] = 10'b1000000101;
    16'b0001001100000000: out_v[61] = 10'b0011100100;
    16'b0001001010001000: out_v[61] = 10'b1110111011;
    16'b0001101010001000: out_v[61] = 10'b1011011011;
    16'b0101011100001000: out_v[61] = 10'b1010000110;
    16'b0001001011001000: out_v[61] = 10'b1110010100;
    16'b0001011100001000: out_v[61] = 10'b1111111101;
    16'b0001011001001000: out_v[61] = 10'b1010111111;
    16'b0000000101001101: out_v[61] = 10'b1011000100;
    16'b0001101011001000: out_v[61] = 10'b1011001010;
    16'b0001101110001000: out_v[61] = 10'b0100101111;
    16'b0101010001000101: out_v[61] = 10'b0010000101;
    16'b0000000101001000: out_v[61] = 10'b1001110111;
    16'b0001000100001000: out_v[61] = 10'b0001001111;
    16'b0101011000000000: out_v[61] = 10'b0111011010;
    16'b0001001110001000: out_v[61] = 10'b0011100011;
    16'b1001001000001000: out_v[61] = 10'b1101010100;
    16'b0001000000001000: out_v[61] = 10'b1011010101;
    16'b0101010000001000: out_v[61] = 10'b1100010101;
    16'b0010001101001101: out_v[61] = 10'b0011101111;
    16'b0000001101001101: out_v[61] = 10'b0110000010;
    16'b0011000101000000: out_v[61] = 10'b0001111101;
    16'b0100011101001101: out_v[61] = 10'b1110011010;
    16'b0110011101000101: out_v[61] = 10'b1101110110;
    16'b0010001001000000: out_v[61] = 10'b1101000111;
    16'b0010001101000101: out_v[61] = 10'b1101100110;
    16'b0010001100001101: out_v[61] = 10'b0011111011;
    16'b0011001101000101: out_v[61] = 10'b0010011101;
    16'b0000001101001000: out_v[61] = 10'b1010111000;
    16'b0010001001000101: out_v[61] = 10'b1010001100;
    16'b0110011001000101: out_v[61] = 10'b0011001111;
    16'b0110011001001101: out_v[61] = 10'b0010011111;
    16'b0010001001001101: out_v[61] = 10'b0110000111;
    16'b0010001101001000: out_v[61] = 10'b1011010010;
    16'b0011001101001101: out_v[61] = 10'b1011101111;
    16'b1100010100001101: out_v[61] = 10'b1000111100;
    16'b0001000101001101: out_v[61] = 10'b0110011000;
    16'b0010001101000000: out_v[61] = 10'b0001100111;
    16'b0000001101000101: out_v[61] = 10'b0101001001;
    16'b0001001111001101: out_v[61] = 10'b1110010111;
    16'b0000001100001101: out_v[61] = 10'b1010001001;
    16'b0000011101001101: out_v[61] = 10'b0110001111;
    16'b0001001100001101: out_v[61] = 10'b0100100100;
    16'b0100010100001101: out_v[61] = 10'b1111111100;
    16'b0000001101001001: out_v[61] = 10'b0011111010;
    16'b0000000100001101: out_v[61] = 10'b0101111010;
    16'b0010001001001000: out_v[61] = 10'b1101100010;
    16'b0110011101001101: out_v[61] = 10'b0011110100;
    16'b0000001101000000: out_v[61] = 10'b0001010110;
    16'b0100011100001101: out_v[61] = 10'b0011110111;
    16'b0000010100001101: out_v[61] = 10'b1010001100;
    16'b0010001101000001: out_v[61] = 10'b0101111111;
    16'b0100011101001000: out_v[61] = 10'b0100111010;
    16'b0100010101001101: out_v[61] = 10'b0110110100;
    16'b0000001100000101: out_v[61] = 10'b1100001001;
    16'b0010011101000101: out_v[61] = 10'b1101111111;
    16'b0000001001000000: out_v[61] = 10'b1010011011;
    16'b0001001001000100: out_v[61] = 10'b1001000011;
    16'b0011101101000000: out_v[61] = 10'b1001001101;
    16'b0001101001001100: out_v[61] = 10'b0000111111;
    16'b0001001011000000: out_v[61] = 10'b0111011101;
    16'b1001001101000000: out_v[61] = 10'b0110000101;
    16'b0001101001000100: out_v[61] = 10'b0111011011;
    16'b0001101101000000: out_v[61] = 10'b0100011011;
    16'b0011001001000000: out_v[61] = 10'b1101000011;
    16'b0001001110000000: out_v[61] = 10'b0011111101;
    16'b0011001101000100: out_v[61] = 10'b0001110011;
    16'b0001001101000001: out_v[61] = 10'b0110110101;
    16'b0001001111000000: out_v[61] = 10'b1111000111;
    16'b0011101111000000: out_v[61] = 10'b0010101011;
    16'b0100011001000000: out_v[61] = 10'b0010111011;
    16'b0000001000000000: out_v[61] = 10'b1110110010;
    16'b0011001110000000: out_v[61] = 10'b0001011011;
    16'b0001001101000000: out_v[61] = 10'b0011000110;
    16'b0011001101000000: out_v[61] = 10'b1101000010;
    16'b0001001010000000: out_v[61] = 10'b0111110010;
    16'b0011001011000000: out_v[61] = 10'b1101010111;
    16'b0001001101000100: out_v[61] = 10'b0110011001;
    16'b0000011001000000: out_v[61] = 10'b0011011111;
    16'b0001101001000000: out_v[61] = 10'b1000111111;
    16'b0011001111000000: out_v[61] = 10'b0111001110;
    16'b0011001100000000: out_v[61] = 10'b1010100010;
    16'b0000001100000000: out_v[61] = 10'b1001111011;
    16'b0001101001001000: out_v[61] = 10'b1000101110;
    16'b0001001011000100: out_v[61] = 10'b0111101011;
    16'b0001101100000000: out_v[61] = 10'b1010011100;
    16'b0011001000000000: out_v[61] = 10'b0010111111;
    16'b0001001001000101: out_v[61] = 10'b0010011011;
    16'b0001101000000000: out_v[61] = 10'b1010101100;
    16'b0001100001001101: out_v[61] = 10'b0100011100;
    16'b0001101101001101: out_v[61] = 10'b1000110011;
    16'b0000001110001101: out_v[61] = 10'b0110110011;
    16'b0001001110001101: out_v[61] = 10'b0011100110;
    16'b0001000111001000: out_v[61] = 10'b0110110010;
    16'b0000001111001000: out_v[61] = 10'b0110001011;
    16'b0001100101001101: out_v[61] = 10'b1010110100;
    16'b0001101001001101: out_v[61] = 10'b1000100001;
    16'b0000101101001000: out_v[61] = 10'b1011011010;
    16'b0001001111001100: out_v[61] = 10'b1110101111;
    16'b0010001111001000: out_v[61] = 10'b1011111110;
    16'b0000100001001101: out_v[61] = 10'b0100110000;
    16'b0001000111001101: out_v[61] = 10'b0111011000;
    16'b0000001101001100: out_v[61] = 10'b1010110111;
    16'b0001101001000101: out_v[61] = 10'b0000110110;
    16'b0010001111000000: out_v[61] = 10'b0111010111;
    16'b0000001111001100: out_v[61] = 10'b1100111111;
    16'b0011000111001000: out_v[61] = 10'b1001011011;
    16'b0000001111001101: out_v[61] = 10'b1111010000;
    16'b0001100001000101: out_v[61] = 10'b1111101000;
    16'b1101011101000000: out_v[61] = 10'b1100011101;
    16'b1101011100000000: out_v[61] = 10'b0110100111;
    16'b0101011100000000: out_v[61] = 10'b1011001010;
    16'b1100011100000000: out_v[61] = 10'b1110010110;
    16'b0000000101000100: out_v[61] = 10'b1011001010;
    16'b0000000100000000: out_v[61] = 10'b1001010111;
    16'b1101011100001000: out_v[61] = 10'b1011111010;
    16'b1101011000000000: out_v[61] = 10'b1011100000;
    16'b0100011101000000: out_v[61] = 10'b1110010011;
    16'b0001000100000000: out_v[61] = 10'b1101011100;
    16'b0000001101000100: out_v[61] = 10'b0111110111;
    16'b0000000101000000: out_v[61] = 10'b1111100111;
    16'b0101011101000100: out_v[61] = 10'b1011100110;
    16'b0001000101000100: out_v[61] = 10'b1111101011;
    16'b0001001011001101: out_v[61] = 10'b1011001011;
    16'b0001011100000000: out_v[61] = 10'b0101011111;
    16'b1101011101001000: out_v[61] = 10'b1110011111;
    16'b0001001000001100: out_v[61] = 10'b0011010111;
    16'b0101011101000000: out_v[61] = 10'b0011001111;
    16'b0001001001001100: out_v[61] = 10'b1001001110;
    16'b0100011100000000: out_v[61] = 10'b0111011110;
    16'b0001101000001101: out_v[61] = 10'b0110000010;
    16'b0000001000000101: out_v[61] = 10'b1011100000;
    16'b0011001100000111: out_v[61] = 10'b0111011100;
    16'b0001000000000000: out_v[61] = 10'b0010111010;
    16'b0000001100000010: out_v[61] = 10'b0010100011;
    16'b0001001000000101: out_v[61] = 10'b1010010110;
    16'b0011001100000101: out_v[61] = 10'b1101000110;
    16'b0001001100000111: out_v[61] = 10'b1101000111;
    16'b0011101100000101: out_v[61] = 10'b0110000111;
    16'b0001101000000100: out_v[61] = 10'b0111111010;
    16'b0011001100000010: out_v[61] = 10'b1100111111;
    16'b0001101000001000: out_v[61] = 10'b1111110011;
    16'b0011001000000101: out_v[61] = 10'b1011000101;
    16'b0011001100000100: out_v[61] = 10'b0111111100;
    16'b0001001100000010: out_v[61] = 10'b0011101110;
    16'b0011001100000110: out_v[61] = 10'b1101111110;
    16'b0011101100000000: out_v[61] = 10'b1101011011;
    16'b0011101000000000: out_v[61] = 10'b0101010011;
    16'b0011001000000100: out_v[61] = 10'b0101111110;
    16'b0001001000000100: out_v[61] = 10'b1001100110;
    16'b0001101000000101: out_v[61] = 10'b1110001111;
    16'b0011000000000000: out_v[61] = 10'b0110010001;
    16'b0011001100000001: out_v[61] = 10'b0111110010;
    16'b0011101100000111: out_v[61] = 10'b0010111110;
    16'b0011101100000100: out_v[61] = 10'b1111011100;
    16'b0001101000001100: out_v[61] = 10'b0010101001;
    16'b0011000101001100: out_v[61] = 10'b0111010111;
    16'b0011100101001100: out_v[61] = 10'b1110110110;
    16'b0011000001000000: out_v[61] = 10'b1000110011;
    16'b0011100101001000: out_v[61] = 10'b0011100011;
    16'b0011101101001100: out_v[61] = 10'b1001100110;
    16'b0011000101001000: out_v[61] = 10'b0010111011;
    16'b0011101111001000: out_v[61] = 10'b0101000001;
    16'b0011001101001100: out_v[61] = 10'b1011111001;
    16'b0011000101001101: out_v[61] = 10'b0011001100;
    16'b0001000101001100: out_v[61] = 10'b0101110000;
    16'b0011101111001101: out_v[61] = 10'b1010110000;
    16'b0011101101001101: out_v[61] = 10'b1101100000;
    16'b0011100101001101: out_v[61] = 10'b1011110000;
    16'b0011101101001000: out_v[61] = 10'b0100101111;
    16'b0011101111001100: out_v[61] = 10'b0111001110;
    16'b0011001101001000: out_v[61] = 10'b0101111010;
    16'b0011100111001000: out_v[61] = 10'b1010011111;
    16'b0001001101000010: out_v[61] = 10'b1010100011;
    16'b0011001101000010: out_v[61] = 10'b1001101111;
    16'b0000001001000101: out_v[61] = 10'b1101011100;
    16'b0011001101000001: out_v[61] = 10'b1101010001;
    16'b0011001001000100: out_v[61] = 10'b0101111111;
    16'b0000001001000001: out_v[61] = 10'b0011101111;
    default: out_v[61] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001000010000010: out_v[62] = 10'b1010011000;
    16'b0000000011000010: out_v[62] = 10'b1000100101;
    16'b0000000010000010: out_v[62] = 10'b0110100001;
    16'b0001000011000010: out_v[62] = 10'b0100100110;
    16'b0000000000000000: out_v[62] = 10'b0111101011;
    16'b0000100010000000: out_v[62] = 10'b0011001101;
    16'b0000000010000000: out_v[62] = 10'b1100011101;
    16'b0001000000000010: out_v[62] = 10'b0001011000;
    16'b0000100011000000: out_v[62] = 10'b0010001100;
    16'b0000000000000010: out_v[62] = 10'b1001001101;
    16'b0000000011000000: out_v[62] = 10'b0011001101;
    16'b0000100011000010: out_v[62] = 10'b1101001110;
    16'b0000100001000000: out_v[62] = 10'b1101100101;
    16'b0000000001000010: out_v[62] = 10'b1100100001;
    16'b0000100000000000: out_v[62] = 10'b1010010101;
    16'b0000000001000000: out_v[62] = 10'b0101111011;
    16'b0000100010000010: out_v[62] = 10'b1011001010;
    16'b0001000001000010: out_v[62] = 10'b1110000100;
    16'b0001100010000010: out_v[62] = 10'b1100110011;
    16'b0001000011000000: out_v[62] = 10'b1101011010;
    16'b0001000000000000: out_v[62] = 10'b1111010000;
    16'b0001000001000000: out_v[62] = 10'b1100110011;
    16'b0000100010001000: out_v[62] = 10'b1010100001;
    16'b0001110011000000: out_v[62] = 10'b1110110101;
    16'b0001100011000000: out_v[62] = 10'b0011111100;
    16'b0001010001000000: out_v[62] = 10'b1011110111;
    16'b0000110011000000: out_v[62] = 10'b1111110011;
    16'b0001100010000000: out_v[62] = 10'b1101100011;
    16'b0001110010000000: out_v[62] = 10'b1001001110;
    16'b0001110001000000: out_v[62] = 10'b0011011011;
    16'b0001100000000000: out_v[62] = 10'b0111110011;
    16'b0001000010000000: out_v[62] = 10'b1100110000;
    16'b0000110000000000: out_v[62] = 10'b1110111101;
    16'b0001110011000010: out_v[62] = 10'b0110011111;
    16'b0001110000000000: out_v[62] = 10'b1011100110;
    16'b0000110010000000: out_v[62] = 10'b0101000011;
    16'b0001100001000000: out_v[62] = 10'b0101001110;
    16'b0001100011000010: out_v[62] = 10'b1110001010;
    16'b0001010000000000: out_v[62] = 10'b0110001010;
    16'b0001000000001000: out_v[62] = 10'b0000110010;
    16'b0001100010001000: out_v[62] = 10'b0110000111;
    16'b0001100001001000: out_v[62] = 10'b1100101111;
    16'b0001100011001000: out_v[62] = 10'b1010111000;
    16'b0001100011010000: out_v[62] = 10'b1100101111;
    16'b0001010010000000: out_v[62] = 10'b1011001100;
    16'b0001110010000010: out_v[62] = 10'b1010101101;
    16'b0001010010000010: out_v[62] = 10'b1011100010;
    16'b0000010010000010: out_v[62] = 10'b0011000011;
    16'b0001000010010000: out_v[62] = 10'b1001100110;
    16'b0000110010000010: out_v[62] = 10'b1111100010;
    16'b0001001010000010: out_v[62] = 10'b0010111001;
    16'b0001001000000010: out_v[62] = 10'b1001100100;
    16'b0001000000001010: out_v[62] = 10'b1000101111;
    default: out_v[62] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1001010100000010: out_v[63] = 10'b1100010101;
    16'b1100010010100000: out_v[63] = 10'b0111101011;
    16'b1100010000000010: out_v[63] = 10'b0001101011;
    16'b0100010100100000: out_v[63] = 10'b1100010111;
    16'b1001010010100000: out_v[63] = 10'b1001001111;
    16'b1001010010100100: out_v[63] = 10'b0111110111;
    16'b1001010010100110: out_v[63] = 10'b0011111011;
    16'b1001010010000010: out_v[63] = 10'b1011001111;
    16'b1100010010000010: out_v[63] = 10'b0101001010;
    16'b1100010100000010: out_v[63] = 10'b0000010111;
    16'b0100010100000010: out_v[63] = 10'b0110010111;
    16'b1001010110100000: out_v[63] = 10'b1110011011;
    16'b1001010000000010: out_v[63] = 10'b1011001000;
    16'b1100010010100110: out_v[63] = 10'b1000111100;
    16'b1000010000000010: out_v[63] = 10'b0101101110;
    16'b1100010010100100: out_v[63] = 10'b1000111011;
    16'b0100010010100000: out_v[63] = 10'b0101111110;
    16'b0001010100000010: out_v[63] = 10'b0010011011;
    16'b0100010100000000: out_v[63] = 10'b0010010111;
    16'b0100010010000010: out_v[63] = 10'b1011111011;
    16'b1100010110100000: out_v[63] = 10'b1101100010;
    16'b0100010010000000: out_v[63] = 10'b1011011001;
    16'b1001000010100010: out_v[63] = 10'b0011110011;
    16'b1001010000100010: out_v[63] = 10'b1011101010;
    16'b0100010000000010: out_v[63] = 10'b1011100000;
    16'b1101010010100110: out_v[63] = 10'b1100101001;
    16'b1001010010100010: out_v[63] = 10'b1011111110;
    16'b0100010110100000: out_v[63] = 10'b0010101110;
    16'b1001010110100110: out_v[63] = 10'b0100001111;
    16'b0100010010100100: out_v[63] = 10'b1011011100;
    16'b0100010000100000: out_v[63] = 10'b1111010001;
    16'b1000010010100000: out_v[63] = 10'b0110111011;
    16'b0000010000000010: out_v[63] = 10'b0001110101;
    16'b1000010100000010: out_v[63] = 10'b1110011111;
    16'b1001010000100000: out_v[63] = 10'b1001100111;
    16'b0100000010100000: out_v[63] = 10'b1011000001;
    16'b1101010000000010: out_v[63] = 10'b0100110110;
    16'b1101010100000010: out_v[63] = 10'b0111010010;
    16'b1001010100100010: out_v[63] = 10'b0000111011;
    16'b0100010000000000: out_v[63] = 10'b0000011010;
    16'b1001010110100010: out_v[63] = 10'b1111111101;
    16'b1001000000000010: out_v[63] = 10'b0100000111;
    16'b0001010100000000: out_v[63] = 10'b0101001101;
    16'b0000000100000000: out_v[63] = 10'b1010000111;
    16'b0000000000000000: out_v[63] = 10'b1100010001;
    16'b0001000000000000: out_v[63] = 10'b1000010111;
    16'b0000010000000000: out_v[63] = 10'b1101110010;
    16'b0000010100000010: out_v[63] = 10'b1010000100;
    16'b0000010100000000: out_v[63] = 10'b0101110111;
    16'b0001010000000000: out_v[63] = 10'b0100011011;
    16'b0101000000000000: out_v[63] = 10'b1100010010;
    16'b0001000100000000: out_v[63] = 10'b0110010100;
    16'b0100000100000000: out_v[63] = 10'b0001001011;
    16'b1100010100000000: out_v[63] = 10'b1101011100;
    16'b1000000100000010: out_v[63] = 10'b1000001010;
    16'b1000010100000000: out_v[63] = 10'b0100011100;
    16'b1000010000100010: out_v[63] = 10'b1111011010;
    16'b1100010000100010: out_v[63] = 10'b0001001100;
    16'b1000010100100010: out_v[63] = 10'b0110110110;
    16'b1100010100100010: out_v[63] = 10'b0000010101;
    16'b0101010000000010: out_v[63] = 10'b0110110100;
    16'b0001010000000010: out_v[63] = 10'b1111011100;
    16'b1100010100010010: out_v[63] = 10'b1101010110;
    16'b0100000000000000: out_v[63] = 10'b0011010101;
    16'b0101010000000000: out_v[63] = 10'b1001110010;
    16'b0100010100100010: out_v[63] = 10'b1110100100;
    16'b0000010100100010: out_v[63] = 10'b1011110111;
    16'b0101010100000010: out_v[63] = 10'b1101010100;
    16'b1100000000000010: out_v[63] = 10'b0011111010;
    16'b1100010000000000: out_v[63] = 10'b0110101011;
    16'b0000010000100010: out_v[63] = 10'b0111001110;
    16'b1100000100000010: out_v[63] = 10'b1000001100;
    16'b1101000000000010: out_v[63] = 10'b1101001000;
    16'b0100010100010000: out_v[63] = 10'b1001001111;
    16'b1000010000100000: out_v[63] = 10'b1110111100;
    16'b1000010000000000: out_v[63] = 10'b0110111110;
    16'b1101000000000000: out_v[63] = 10'b1100001011;
    16'b1001000000000000: out_v[63] = 10'b0111011100;
    16'b1001010000000000: out_v[63] = 10'b1000101110;
    16'b1001000100000000: out_v[63] = 10'b0010110101;
    16'b0100000100000010: out_v[63] = 10'b0011001111;
    16'b1101010100000000: out_v[63] = 10'b1011100110;
    16'b1101010100010000: out_v[63] = 10'b1011101011;
    16'b1100000100000000: out_v[63] = 10'b0011010010;
    16'b1101010000000000: out_v[63] = 10'b0000111011;
    16'b1000000100000000: out_v[63] = 10'b1101001000;
    16'b0101000000010000: out_v[63] = 10'b1100011101;
    16'b1101000000010000: out_v[63] = 10'b1100010010;
    16'b0101010000010000: out_v[63] = 10'b1000011000;
    16'b1001010100100000: out_v[63] = 10'b0001001110;
    16'b0101000000000010: out_v[63] = 10'b0111001100;
    16'b1101000100000000: out_v[63] = 10'b1100000101;
    16'b0101010100000000: out_v[63] = 10'b1011111000;
    16'b1100001100000000: out_v[63] = 10'b1111110010;
    16'b1100000100010000: out_v[63] = 10'b1110000000;
    16'b1001010100000000: out_v[63] = 10'b0010101110;
    16'b1101010100100000: out_v[63] = 10'b0111101100;
    16'b1101001100000000: out_v[63] = 10'b0100011110;
    16'b1101000100000010: out_v[63] = 10'b0011111111;
    16'b1100000000000000: out_v[63] = 10'b0110110001;
    16'b1101000100010000: out_v[63] = 10'b1010100111;
    16'b0101000100000000: out_v[63] = 10'b1101100100;
    16'b0001000100100010: out_v[63] = 10'b0011110011;
    16'b0001000000000010: out_v[63] = 10'b0000010011;
    16'b0001000100000010: out_v[63] = 10'b0110101000;
    16'b0000000000000010: out_v[63] = 10'b0010110001;
    16'b1100000100001010: out_v[63] = 10'b0100110010;
    16'b0000000100000010: out_v[63] = 10'b1000110001;
    16'b1100000100100010: out_v[63] = 10'b1001100110;
    16'b1000000100010010: out_v[63] = 10'b0011011111;
    16'b1000000000000010: out_v[63] = 10'b1100111010;
    16'b1000000100100010: out_v[63] = 10'b0001100101;
    16'b1001000100000010: out_v[63] = 10'b0110011000;
    16'b1000000000100010: out_v[63] = 10'b0000101110;
    16'b0000000100100010: out_v[63] = 10'b1000000111;
    16'b1001000100100010: out_v[63] = 10'b0100011000;
    16'b0100000000000010: out_v[63] = 10'b0011100011;
    16'b1001000000100010: out_v[63] = 10'b1000111110;
    16'b1000000000000000: out_v[63] = 10'b0111000101;
    16'b1100000000100010: out_v[63] = 10'b0011111101;
    16'b0001010110000100: out_v[63] = 10'b0011001110;
    16'b0001010000100000: out_v[63] = 10'b1001110000;
    16'b1001000110000000: out_v[63] = 10'b0010011000;
    16'b1100000100001000: out_v[63] = 10'b0111001111;
    16'b1101000100001000: out_v[63] = 10'b1100100111;
    16'b1000000100001000: out_v[63] = 10'b0000110111;
    16'b0100000100010000: out_v[63] = 10'b1011010100;
    16'b1100000100011000: out_v[63] = 10'b1101111011;
    16'b1001000100001000: out_v[63] = 10'b0110101011;
    16'b1001000100010000: out_v[63] = 10'b1000110010;
    16'b0001010010000110: out_v[63] = 10'b0110101000;
    16'b0000000100001010: out_v[63] = 10'b1011101111;
    16'b1000000100001010: out_v[63] = 10'b0100111101;
    16'b1100000000001000: out_v[63] = 10'b0111000011;
    16'b0100000000001000: out_v[63] = 10'b1100101100;
    16'b0100000100001000: out_v[63] = 10'b0001010110;
    16'b1100000000001010: out_v[63] = 10'b0001100010;
    16'b0100000100001010: out_v[63] = 10'b0011001010;
    16'b1000000000001010: out_v[63] = 10'b1111010011;
    16'b1001000100001010: out_v[63] = 10'b1111000010;
    default: out_v[63] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100010110010000: out_v[64] = 10'b0011011100;
    16'b0100010111000100: out_v[64] = 10'b1010010110;
    16'b0000010000000100: out_v[64] = 10'b1101100010;
    16'b0100100111001100: out_v[64] = 10'b0010111001;
    16'b0100000111000100: out_v[64] = 10'b0110011011;
    16'b0110000111000100: out_v[64] = 10'b1010101111;
    16'b0110000111000000: out_v[64] = 10'b1110010111;
    16'b0100010111010000: out_v[64] = 10'b1000111101;
    16'b0100010110000100: out_v[64] = 10'b1111100001;
    16'b0000110110000100: out_v[64] = 10'b1100101110;
    16'b0000010001000100: out_v[64] = 10'b0111000111;
    16'b0100110111001100: out_v[64] = 10'b1111110111;
    16'b0000010011000100: out_v[64] = 10'b1011010111;
    16'b0100110110001100: out_v[64] = 10'b0110011010;
    16'b0110010111000100: out_v[64] = 10'b1111100110;
    16'b0000010110000100: out_v[64] = 10'b1111111011;
    16'b0100010111010100: out_v[64] = 10'b0011110011;
    16'b0100010011000100: out_v[64] = 10'b0011001111;
    16'b0110100111001100: out_v[64] = 10'b1100111111;
    16'b0110110111001100: out_v[64] = 10'b1010010111;
    16'b0000010111000100: out_v[64] = 10'b1001110100;
    16'b0100000111001100: out_v[64] = 10'b1111001011;
    16'b0110010111000000: out_v[64] = 10'b1100111001;
    16'b0100000101000100: out_v[64] = 10'b1110110011;
    16'b0100110110000100: out_v[64] = 10'b1011010101;
    16'b0000110000000100: out_v[64] = 10'b1000111111;
    16'b0000010001010000: out_v[64] = 10'b1000110101;
    16'b0000110000001100: out_v[64] = 10'b1001100001;
    16'b0100010110000000: out_v[64] = 10'b1011001001;
    16'b0100010111000000: out_v[64] = 10'b0000100101;
    16'b0110110110001100: out_v[64] = 10'b0001100101;
    16'b0100010111001100: out_v[64] = 10'b0010111101;
    16'b0000010100000100: out_v[64] = 10'b1111111101;
    16'b0000010010000100: out_v[64] = 10'b1000011111;
    16'b0100110111000100: out_v[64] = 10'b1101110100;
    16'b0000110100001100: out_v[64] = 10'b0011011111;
    16'b0100010100100000: out_v[64] = 10'b0010010010;
    16'b0100000110100000: out_v[64] = 10'b0010101011;
    16'b0100000010100000: out_v[64] = 10'b1000001011;
    16'b0100010110100000: out_v[64] = 10'b0011100010;
    16'b0100000100100000: out_v[64] = 10'b1010110101;
    16'b0100000011100000: out_v[64] = 10'b0011011011;
    16'b0100000010000000: out_v[64] = 10'b1110001100;
    16'b0100000000100000: out_v[64] = 10'b0110101010;
    16'b0000000000100000: out_v[64] = 10'b1001011010;
    16'b0100010010100000: out_v[64] = 10'b1100000001;
    16'b0000000011100000: out_v[64] = 10'b1011001110;
    16'b0000000001100000: out_v[64] = 10'b0001000111;
    16'b0100000111100000: out_v[64] = 10'b1101010001;
    16'b0000010000100000: out_v[64] = 10'b0011111100;
    16'b0100010111100000: out_v[64] = 10'b0001101100;
    16'b0100000011000000: out_v[64] = 10'b0110111111;
    16'b0000000010100000: out_v[64] = 10'b0010011011;
    16'b0001000000100000: out_v[64] = 10'b1110100011;
    16'b0100010000100000: out_v[64] = 10'b1100100001;
    16'b0000010100100000: out_v[64] = 10'b0011111111;
    16'b0100100111100000: out_v[64] = 10'b1010100001;
    16'b0100100101100000: out_v[64] = 10'b0101111011;
    16'b0000100101100000: out_v[64] = 10'b1010111111;
    16'b0000100101110000: out_v[64] = 10'b1111001010;
    16'b0000000101110000: out_v[64] = 10'b1010101110;
    16'b0000000000110000: out_v[64] = 10'b0101110111;
    16'b0000010001110000: out_v[64] = 10'b1010001000;
    16'b0000000001110000: out_v[64] = 10'b0010011011;
    16'b0100110111110000: out_v[64] = 10'b1001111111;
    16'b0000000001100100: out_v[64] = 10'b0101001110;
    16'b0100100111110000: out_v[64] = 10'b0100010110;
    16'b0100110111100000: out_v[64] = 10'b1011101101;
    16'b0100000101110000: out_v[64] = 10'b0001111100;
    16'b0000100001110000: out_v[64] = 10'b1001100011;
    16'b0100000110110000: out_v[64] = 10'b1111100100;
    16'b0000100000110000: out_v[64] = 10'b1111001111;
    16'b0000000101100000: out_v[64] = 10'b1101001110;
    16'b0100010111110000: out_v[64] = 10'b1011001110;
    16'b0000000001010000: out_v[64] = 10'b0101011110;
    16'b0000000001110100: out_v[64] = 10'b0110110011;
    16'b0000100001100000: out_v[64] = 10'b0011000010;
    16'b0100000111110000: out_v[64] = 10'b1101001000;
    16'b0000000000110100: out_v[64] = 10'b1010000110;
    16'b0000000011110000: out_v[64] = 10'b0110011011;
    16'b0100000101100000: out_v[64] = 10'b0101010100;
    16'b0000000100110000: out_v[64] = 10'b1111111011;
    16'b0000100000100000: out_v[64] = 10'b0001011101;
    16'b0000010000110000: out_v[64] = 10'b0100111010;
    16'b0100100110100000: out_v[64] = 10'b0100101101;
    16'b0100100100100000: out_v[64] = 10'b1000100001;
    16'b0100100011100000: out_v[64] = 10'b1000111011;
    16'b0000000100100000: out_v[64] = 10'b1010001101;
    16'b0100100110110000: out_v[64] = 10'b0110101110;
    16'b0000100001100100: out_v[64] = 10'b1110000011;
    16'b0000010101110000: out_v[64] = 10'b1001000110;
    16'b0100000110110100: out_v[64] = 10'b1001100110;
    16'b0100010100010000: out_v[64] = 10'b1100011010;
    16'b0100010100000000: out_v[64] = 10'b1100001111;
    16'b0000010111010000: out_v[64] = 10'b1111110011;
    16'b0000010000010000: out_v[64] = 10'b0101110000;
    16'b0000010000000000: out_v[64] = 10'b0110110001;
    16'b0100010101010000: out_v[64] = 10'b1010001011;
    16'b0100110110010000: out_v[64] = 10'b1101011100;
    16'b0000010001000000: out_v[64] = 10'b0011110010;
    16'b0100110100000000: out_v[64] = 10'b0111011100;
    16'b0100110110000000: out_v[64] = 10'b0111011010;
    16'b0100010101000000: out_v[64] = 10'b1000001100;
    16'b0100110110100000: out_v[64] = 10'b1010111010;
    16'b0000110000010000: out_v[64] = 10'b1000110110;
    16'b0000010111110000: out_v[64] = 10'b1011101011;
    16'b0100000111010000: out_v[64] = 10'b0110001111;
    16'b0100000101000000: out_v[64] = 10'b0000110011;
    16'b0100110100010000: out_v[64] = 10'b1101011011;
    16'b0100010001010000: out_v[64] = 10'b0111100001;
    16'b0000010011010000: out_v[64] = 10'b1001110110;
    16'b0100010101100000: out_v[64] = 10'b1100001101;
    16'b0100010000010000: out_v[64] = 10'b1111101010;
    16'b0000010100000000: out_v[64] = 10'b1001100111;
    16'b0100010010010000: out_v[64] = 10'b1110100100;
    16'b0100000101010000: out_v[64] = 10'b0111001100;
    16'b0000010001100000: out_v[64] = 10'b0001101011;
    16'b0100010000000000: out_v[64] = 10'b1001101110;
    16'b0000010101100000: out_v[64] = 10'b0101110011;
    16'b0000010111100000: out_v[64] = 10'b0100111101;
    16'b0100010001000000: out_v[64] = 10'b0110011111;
    16'b0000010101000000: out_v[64] = 10'b1100110001;
    16'b0100010010000000: out_v[64] = 10'b1101001100;
    16'b0000000001000000: out_v[64] = 10'b1001100010;
    16'b0100010110110000: out_v[64] = 10'b1111101110;
    16'b0000000000010000: out_v[64] = 10'b0011110110;
    16'b0000010001110100: out_v[64] = 10'b1111101001;
    16'b0000000000111000: out_v[64] = 10'b0011100111;
    16'b0000010010110000: out_v[64] = 10'b1001100110;
    16'b0000000001111000: out_v[64] = 10'b1011001111;
    16'b0000000000000000: out_v[64] = 10'b1000111111;
    16'b0100000101111000: out_v[64] = 10'b0010011110;
    16'b0000000100111000: out_v[64] = 10'b0011010111;
    16'b0000000001011000: out_v[64] = 10'b0010110001;
    16'b0000000001111100: out_v[64] = 10'b0110110001;
    16'b0100010010110000: out_v[64] = 10'b0111111100;
    16'b0000010000110100: out_v[64] = 10'b0110000000;
    16'b0000000000111100: out_v[64] = 10'b0011101010;
    16'b0000000000100100: out_v[64] = 10'b0010110000;
    16'b0000010010100000: out_v[64] = 10'b0101010000;
    16'b0100000011110000: out_v[64] = 10'b0001110010;
    16'b0100000000000000: out_v[64] = 10'b0010111000;
    16'b0100000001000000: out_v[64] = 10'b1000101010;
    16'b0100000110000000: out_v[64] = 10'b1010101100;
    16'b0100000111000000: out_v[64] = 10'b0111110010;
    16'b0100000001100000: out_v[64] = 10'b1111000101;
    16'b0000010110000000: out_v[64] = 10'b1011100101;
    16'b0000010110100000: out_v[64] = 10'b0111100001;
    16'b0000010111000000: out_v[64] = 10'b0011110010;
    16'b0000010011000000: out_v[64] = 10'b0011001111;
    16'b0000110000000000: out_v[64] = 10'b1010100101;
    16'b0000010010000000: out_v[64] = 10'b1010011011;
    16'b0000010011100000: out_v[64] = 10'b0110101010;
    16'b0000010010010000: out_v[64] = 10'b1001001110;
    16'b0000110000011000: out_v[64] = 10'b1001110111;
    16'b0100000100000000: out_v[64] = 10'b1001011100;
    16'b0101000111100000: out_v[64] = 10'b1101000110;
    16'b0010100001111100: out_v[64] = 10'b0111001110;
    16'b0100000011110100: out_v[64] = 10'b1100101011;
    16'b0000000011000000: out_v[64] = 10'b1100110010;
    16'b0000100001110100: out_v[64] = 10'b0110010011;
    16'b0000000010110000: out_v[64] = 10'b0001011111;
    16'b0000000011110100: out_v[64] = 10'b0100111001;
    16'b0000000001010100: out_v[64] = 10'b0101101010;
    16'b0100000111110100: out_v[64] = 10'b1001001000;
    16'b0000000011010000: out_v[64] = 10'b1100011000;
    16'b0000000001000100: out_v[64] = 10'b1110011100;
    16'b0100000011010000: out_v[64] = 10'b1111100010;
    16'b0000100001010000: out_v[64] = 10'b1110010101;
    16'b0010000001110100: out_v[64] = 10'b1010101011;
    16'b0100010110011000: out_v[64] = 10'b0101000110;
    16'b0100010111011000: out_v[64] = 10'b0111011010;
    16'b0100000110011000: out_v[64] = 10'b0111010001;
    16'b0100000111011000: out_v[64] = 10'b0111010010;
    16'b0100000001010000: out_v[64] = 10'b0110100111;
    16'b0100010110010100: out_v[64] = 10'b0001111111;
    16'b0100000110010000: out_v[64] = 10'b1011111001;
    16'b0100010111011100: out_v[64] = 10'b0101000111;
    16'b0100000111001000: out_v[64] = 10'b1011010110;
    16'b0100000001011000: out_v[64] = 10'b1001111101;
    16'b0100010110110100: out_v[64] = 10'b0100001100;
    16'b0100000111011100: out_v[64] = 10'b0110111010;
    16'b0100000111111000: out_v[64] = 10'b0111001101;
    16'b0100010110111000: out_v[64] = 10'b0111111111;
    16'b0100010111110100: out_v[64] = 10'b1110001000;
    16'b0000010011110100: out_v[64] = 10'b0111101111;
    16'b0100010011100000: out_v[64] = 10'b1100110101;
    16'b0000010010110100: out_v[64] = 10'b0000011100;
    16'b0000010110110000: out_v[64] = 10'b1101100110;
    16'b0000010111110100: out_v[64] = 10'b0011011001;
    16'b0000010011110000: out_v[64] = 10'b0100110111;
    16'b0100000111111100: out_v[64] = 10'b1101100111;
    16'b0000000111010000: out_v[64] = 10'b1001101101;
    16'b0000000111000000: out_v[64] = 10'b1110101000;
    16'b0000000111100000: out_v[64] = 10'b0001110111;
    16'b0000010110010000: out_v[64] = 10'b1100000110;
    16'b0000000111111000: out_v[64] = 10'b1011110011;
    16'b0000000111110000: out_v[64] = 10'b1111000000;
    16'b0100010111111100: out_v[64] = 10'b1110000000;
    16'b0100000110111000: out_v[64] = 10'b1000001011;
    16'b0100000110111100: out_v[64] = 10'b1001100111;
    default: out_v[64] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000010000101100: out_v[65] = 10'b1000011001;
    16'b0000011000011111: out_v[65] = 10'b1101111111;
    16'b0000010000101011: out_v[65] = 10'b1111000111;
    16'b0000010000001101: out_v[65] = 10'b0010011011;
    16'b0000010000101101: out_v[65] = 10'b1111011100;
    16'b1100010001011111: out_v[65] = 10'b0011111110;
    16'b1100010001010111: out_v[65] = 10'b1001100111;
    16'b1100011001011111: out_v[65] = 10'b1011010110;
    16'b0000010000111111: out_v[65] = 10'b0110001001;
    16'b0000010000111011: out_v[65] = 10'b1110100011;
    16'b1100010001111111: out_v[65] = 10'b1111101010;
    16'b0000010000011111: out_v[65] = 10'b0100001111;
    16'b0000010001011111: out_v[65] = 10'b0110010011;
    16'b1100010000011111: out_v[65] = 10'b0011111101;
    16'b0000010000101111: out_v[65] = 10'b1000101011;
    16'b1100010001011011: out_v[65] = 10'b0111101011;
    16'b0000010000001111: out_v[65] = 10'b1001101001;
    16'b0000000000011111: out_v[65] = 10'b0001011100;
    16'b0000000000000100: out_v[65] = 10'b1011001001;
    16'b0000010000011011: out_v[65] = 10'b0001001111;
    16'b0000000000101011: out_v[65] = 10'b1100101111;
    16'b1100011001010111: out_v[65] = 10'b1111000110;
    16'b1100001001011111: out_v[65] = 10'b0000111101;
    16'b0000010000001011: out_v[65] = 10'b1100100001;
    16'b1100001001010111: out_v[65] = 10'b1011111011;
    16'b0000000000111011: out_v[65] = 10'b0100001100;
    16'b0000010000101001: out_v[65] = 10'b1000100011;
    16'b0000000000001100: out_v[65] = 10'b1001011111;
    16'b1110010001011111: out_v[65] = 10'b1011011111;
    16'b1100010000111011: out_v[65] = 10'b1010101111;
    16'b1100000001011111: out_v[65] = 10'b1110010011;
    16'b1100011001111111: out_v[65] = 10'b1111101011;
    16'b0000010000001100: out_v[65] = 10'b0010010010;
    16'b1110010001111111: out_v[65] = 10'b1100111010;
    16'b1100010001111011: out_v[65] = 10'b1110010010;
    16'b1100011001011101: out_v[65] = 10'b0101101110;
    16'b0000010000101000: out_v[65] = 10'b0100101011;
    16'b1100010000111111: out_v[65] = 10'b0111100100;
    16'b0000000000101111: out_v[65] = 10'b1110010101;
    16'b0000000000000000: out_v[65] = 10'b0001111010;
    16'b0000000000101000: out_v[65] = 10'b1010101000;
    16'b0000000000101100: out_v[65] = 10'b0000001110;
    16'b0000000000100100: out_v[65] = 10'b1111100001;
    16'b0000010000000100: out_v[65] = 10'b1011001010;
    16'b0000000000010000: out_v[65] = 10'b0000111011;
    16'b0000000000001000: out_v[65] = 10'b1011100100;
    16'b0000001000010000: out_v[65] = 10'b1000101011;
    16'b0000000000100000: out_v[65] = 10'b0001111100;
    16'b0000000000001001: out_v[65] = 10'b1000101011;
    16'b0000010000001000: out_v[65] = 10'b1001100111;
    16'b0000010010001000: out_v[65] = 10'b1100100101;
    16'b0000010000000000: out_v[65] = 10'b0010110100;
    16'b0000000010001000: out_v[65] = 10'b0100010100;
    16'b0000000001011010: out_v[65] = 10'b1011010110;
    16'b0000010000001001: out_v[65] = 10'b1011000001;
    16'b0000010001011000: out_v[65] = 10'b1011111100;
    16'b0000010000011000: out_v[65] = 10'b1100100111;
    16'b0000010010001100: out_v[65] = 10'b1110010100;
    16'b0000000010001001: out_v[65] = 10'b0101100101;
    16'b0000000001001000: out_v[65] = 10'b1011010011;
    16'b0000000000000001: out_v[65] = 10'b0000111101;
    16'b0000010001001000: out_v[65] = 10'b1110110011;
    16'b0000010010000000: out_v[65] = 10'b1011100101;
    16'b0000010001011010: out_v[65] = 10'b0111111110;
    16'b0000000001000000: out_v[65] = 10'b1100011001;
    16'b1100000001011010: out_v[65] = 10'b0110111011;
    16'b0000000010000000: out_v[65] = 10'b1110111110;
    16'b1100010001011010: out_v[65] = 10'b0111100001;
    16'b0000010001000000: out_v[65] = 10'b1101110111;
    16'b0000000001011000: out_v[65] = 10'b0101010011;
    16'b1100010001011000: out_v[65] = 10'b0011110110;
    16'b1100000001010011: out_v[65] = 10'b1010111001;
    16'b0000010000000001: out_v[65] = 10'b0000111100;
    16'b0000000010001100: out_v[65] = 10'b0100000110;
    16'b0000010001101000: out_v[65] = 10'b1110000011;
    16'b0000010001001100: out_v[65] = 10'b0011011101;
    16'b0000000000101001: out_v[65] = 10'b1101000011;
    16'b0000010001011100: out_v[65] = 10'b1010010011;
    16'b0000000000011000: out_v[65] = 10'b1111001001;
    16'b0000010000111000: out_v[65] = 10'b1011001011;
    16'b0000000000101101: out_v[65] = 10'b0110001011;
    16'b0000010000111001: out_v[65] = 10'b1101011010;
    16'b0000010000100000: out_v[65] = 10'b1001110011;
    16'b0000010001111000: out_v[65] = 10'b1110000011;
    16'b0000010001000100: out_v[65] = 10'b1011011111;
    16'b0000010001101100: out_v[65] = 10'b0101101111;
    16'b0000010000100100: out_v[65] = 10'b1110010000;
    16'b0000010000100101: out_v[65] = 10'b1101100111;
    16'b0000001000011001: out_v[65] = 10'b1000111010;
    16'b0000000000011101: out_v[65] = 10'b0001111011;
    16'b0000001000011111: out_v[65] = 10'b0000011000;
    16'b0000000000011001: out_v[65] = 10'b0001100010;
    16'b0000010000110001: out_v[65] = 10'b1011001001;
    16'b0000000000000101: out_v[65] = 10'b1110001101;
    16'b0000001000010001: out_v[65] = 10'b0001111001;
    16'b0000000000000011: out_v[65] = 10'b0010111011;
    16'b0000010000000011: out_v[65] = 10'b0111001001;
    16'b0000010000110011: out_v[65] = 10'b1001011111;
    16'b0000010000100001: out_v[65] = 10'b0100011101;
    16'b0000010000010001: out_v[65] = 10'b0111111000;
    16'b0000010000010011: out_v[65] = 10'b0011000101;
    16'b0000001000011101: out_v[65] = 10'b0011110110;
    16'b0000000000100001: out_v[65] = 10'b0100010111;
    16'b0000000000010001: out_v[65] = 10'b0110011100;
    16'b0000001000010101: out_v[65] = 10'b1001001111;
    16'b0000001000010011: out_v[65] = 10'b1001011111;
    16'b0000000000010011: out_v[65] = 10'b0011011010;
    16'b0000000000100101: out_v[65] = 10'b1101000110;
    16'b0000000000001101: out_v[65] = 10'b0010000111;
    16'b0000000000110001: out_v[65] = 10'b1001111111;
    16'b0000011000110011: out_v[65] = 10'b1011011101;
    16'b0000000000010101: out_v[65] = 10'b1100001001;
    16'b1100000000000001: out_v[65] = 10'b1011101110;
    16'b0000000000111001: out_v[65] = 10'b0111110011;
    16'b0000001000011011: out_v[65] = 10'b0011110111;
    16'b0000001000010100: out_v[65] = 10'b0100011101;
    16'b0000011000111101: out_v[65] = 10'b0000100110;
    16'b0000010000111101: out_v[65] = 10'b1001100100;
    16'b0000011000011101: out_v[65] = 10'b0110111110;
    16'b0000011000010101: out_v[65] = 10'b0101110010;
    16'b0000011000111100: out_v[65] = 10'b1110010010;
    16'b0000011000111001: out_v[65] = 10'b1111111010;
    16'b0000010000111100: out_v[65] = 10'b0001110110;
    16'b0000000000010100: out_v[65] = 10'b0100110101;
    16'b0000001001011100: out_v[65] = 10'b1111010101;
    16'b0000001001010100: out_v[65] = 10'b1011110100;
    16'b0000011000011100: out_v[65] = 10'b1111110110;
    16'b0000001000011100: out_v[65] = 10'b0100101010;
    16'b0000001000111101: out_v[65] = 10'b1110100010;
    16'b0000011000101001: out_v[65] = 10'b0001101101;
    16'b1100001000010100: out_v[65] = 10'b0111100010;
    16'b0000010000001010: out_v[65] = 10'b1001011010;
    16'b0000010000000101: out_v[65] = 10'b0110011100;
    16'b0000010000001110: out_v[65] = 10'b1111110010;
    16'b0000010000000010: out_v[65] = 10'b0111110001;
    16'b0000000000001111: out_v[65] = 10'b1001111110;
    16'b0000000000001011: out_v[65] = 10'b1001101011;
    16'b0000010000000111: out_v[65] = 10'b1101011010;
    16'b0000000000001110: out_v[65] = 10'b0100111111;
    16'b0000010010000011: out_v[65] = 10'b1111100011;
    16'b0000010000100110: out_v[65] = 10'b1111110011;
    16'b0000000000011100: out_v[65] = 10'b0100010101;
    16'b0000100000011110: out_v[65] = 10'b1100111110;
    16'b0000000000111100: out_v[65] = 10'b1111010000;
    16'b0000010000101110: out_v[65] = 10'b0101100010;
    16'b0000000000010110: out_v[65] = 10'b1110101001;
    16'b0000000000001010: out_v[65] = 10'b0110100010;
    16'b0000000000011010: out_v[65] = 10'b1111000001;
    16'b0000000000000110: out_v[65] = 10'b0010001100;
    16'b0000000000011110: out_v[65] = 10'b0011101111;
    16'b0000010000110110: out_v[65] = 10'b1010110000;
    16'b0000011000111000: out_v[65] = 10'b1000001011;
    16'b0000010000111110: out_v[65] = 10'b1100010011;
    16'b0000010000101010: out_v[65] = 10'b1000101110;
    16'b0000000000111000: out_v[65] = 10'b0011010111;
    16'b0000000000111010: out_v[65] = 10'b0111011001;
    16'b0000001000011000: out_v[65] = 10'b0011100010;
    16'b0000001000111000: out_v[65] = 10'b1100001111;
    16'b0000010000011100: out_v[65] = 10'b0101110010;
    16'b0000001000111100: out_v[65] = 10'b1100110010;
    16'b0000010000111010: out_v[65] = 10'b1001011011;
    16'b0000001000011110: out_v[65] = 10'b1101011010;
    16'b0000000000101010: out_v[65] = 10'b0100001101;
    16'b0000001001011110: out_v[65] = 10'b0101010011;
    16'b0000000000011011: out_v[65] = 10'b1001000011;
    16'b0000000000010111: out_v[65] = 10'b0111101110;
    default: out_v[65] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000100000100000: out_v[66] = 10'b1001101011;
    16'b0001100000000010: out_v[66] = 10'b1000010011;
    16'b0001110000100010: out_v[66] = 10'b0101000001;
    16'b0000110000000010: out_v[66] = 10'b1010110111;
    16'b0000110000100000: out_v[66] = 10'b1001011001;
    16'b0000010000100010: out_v[66] = 10'b1111100010;
    16'b0001100000100010: out_v[66] = 10'b1000011101;
    16'b0001010000000010: out_v[66] = 10'b1111010011;
    16'b0000010000000000: out_v[66] = 10'b1010001001;
    16'b0001110000000010: out_v[66] = 10'b1010010110;
    16'b0000100000000010: out_v[66] = 10'b0011110111;
    16'b0000010000100000: out_v[66] = 10'b0100010110;
    16'b0000000000000010: out_v[66] = 10'b0010011011;
    16'b0000100000000000: out_v[66] = 10'b0110010111;
    16'b0000111000000010: out_v[66] = 10'b0110110100;
    16'b0000111000100010: out_v[66] = 10'b0001001001;
    16'b0000110000000000: out_v[66] = 10'b1010101001;
    16'b0000010000000010: out_v[66] = 10'b1000110110;
    16'b0000110000100010: out_v[66] = 10'b1001000011;
    16'b0000011000000010: out_v[66] = 10'b0011110100;
    16'b0000111000100000: out_v[66] = 10'b1101000110;
    16'b0001111000100010: out_v[66] = 10'b1010010111;
    16'b0001000000000010: out_v[66] = 10'b0001001111;
    16'b0001010000100010: out_v[66] = 10'b0110000011;
    16'b0000000000100000: out_v[66] = 10'b1101000101;
    16'b0001000000100010: out_v[66] = 10'b1101000011;
    16'b0000100000100010: out_v[66] = 10'b0101001000;
    16'b0001111000000010: out_v[66] = 10'b0011101011;
    16'b0000011000100010: out_v[66] = 10'b0101011100;
    16'b0000000000000000: out_v[66] = 10'b1000101010;
    16'b0001000000100000: out_v[66] = 10'b1010101100;
    16'b0000001000100000: out_v[66] = 10'b0101001010;
    16'b0000101000100000: out_v[66] = 10'b1101100010;
    16'b0000011000000000: out_v[66] = 10'b1001101010;
    16'b0000001000000000: out_v[66] = 10'b1100011110;
    16'b0000011000100000: out_v[66] = 10'b0110110100;
    16'b0000101000000000: out_v[66] = 10'b1101010110;
    16'b0000000000100010: out_v[66] = 10'b0101010100;
    16'b0001100000100000: out_v[66] = 10'b1001111100;
    16'b0000111000000000: out_v[66] = 10'b1110001000;
    16'b0001000000000000: out_v[66] = 10'b0001110000;
    16'b0000001000000010: out_v[66] = 10'b0001011101;
    16'b0001010000000000: out_v[66] = 10'b0011110011;
    16'b0001100000000000: out_v[66] = 10'b1110100010;
    16'b0001110000100000: out_v[66] = 10'b1101010010;
    16'b0001110000000000: out_v[66] = 10'b0000111011;
    16'b0001010000100000: out_v[66] = 10'b0110000110;
    16'b0001011000000000: out_v[66] = 10'b0010111000;
    16'b0010010000000000: out_v[66] = 10'b0111000000;
    default: out_v[66] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000110110010000: out_v[67] = 10'b1000110011;
    16'b0000110100000110: out_v[67] = 10'b1111010011;
    16'b0010110100010110: out_v[67] = 10'b1010100011;
    16'b0000110100010110: out_v[67] = 10'b0010000001;
    16'b0000110100010010: out_v[67] = 10'b1110011100;
    16'b0001110110000000: out_v[67] = 10'b0011100011;
    16'b0001110010000110: out_v[67] = 10'b0000110000;
    16'b0000110100010100: out_v[67] = 10'b1010001111;
    16'b0000000000000110: out_v[67] = 10'b0101000110;
    16'b0000000100010100: out_v[67] = 10'b1101001110;
    16'b0001110010000000: out_v[67] = 10'b1101000011;
    16'b0010110100000110: out_v[67] = 10'b1101000001;
    16'b0011110110010000: out_v[67] = 10'b1011001101;
    16'b0010110110010110: out_v[67] = 10'b1011011011;
    16'b0000110010000000: out_v[67] = 10'b1101100011;
    16'b0000000100010110: out_v[67] = 10'b1000000111;
    16'b0000110110000010: out_v[67] = 10'b1100001010;
    16'b0000110110010110: out_v[67] = 10'b1111001010;
    16'b0000110010000110: out_v[67] = 10'b1111001000;
    16'b0000110000000110: out_v[67] = 10'b0110000111;
    16'b0001010010000000: out_v[67] = 10'b1101010010;
    16'b0000000110010000: out_v[67] = 10'b1001111100;
    16'b0000000000010110: out_v[67] = 10'b0011010111;
    16'b0000010100010110: out_v[67] = 10'b1011100110;
    16'b0000110100000100: out_v[67] = 10'b1110111111;
    16'b0000110110000000: out_v[67] = 10'b0100001011;
    16'b0000110110000110: out_v[67] = 10'b0111110010;
    16'b0001010010000110: out_v[67] = 10'b0110011011;
    16'b0000110110010010: out_v[67] = 10'b1100001001;
    16'b0001110010000010: out_v[67] = 10'b0011001110;
    16'b0000000100010000: out_v[67] = 10'b0001100111;
    16'b0001110110000110: out_v[67] = 10'b1011011101;
    16'b0000000100010010: out_v[67] = 10'b1000100110;
    16'b0001010000000000: out_v[67] = 10'b1000110000;
    16'b0010110110010000: out_v[67] = 10'b0000011011;
    16'b0000110100010000: out_v[67] = 10'b1101100010;
    16'b0001110110010000: out_v[67] = 10'b1001110110;
    16'b0011110010000110: out_v[67] = 10'b1110001000;
    16'b0000100100010110: out_v[67] = 10'b1011000110;
    16'b0011010010000110: out_v[67] = 10'b1011000011;
    16'b0000010010000000: out_v[67] = 10'b0101001011;
    16'b0010000100010110: out_v[67] = 10'b1001000011;
    16'b0001010010000010: out_v[67] = 10'b1010110001;
    16'b0011110110010110: out_v[67] = 10'b0100101011;
    16'b0001110110010110: out_v[67] = 10'b0110010011;
    16'b0010000000000000: out_v[67] = 10'b1000001010;
    16'b0000000000000000: out_v[67] = 10'b0111100000;
    16'b0011000000000000: out_v[67] = 10'b0111110010;
    16'b0010010000000000: out_v[67] = 10'b0100011100;
    16'b0000010000000000: out_v[67] = 10'b0100101110;
    16'b0010000100010000: out_v[67] = 10'b0010010111;
    16'b0001000010000000: out_v[67] = 10'b0010110100;
    16'b0011000100010000: out_v[67] = 10'b0011001001;
    16'b0001000000010000: out_v[67] = 10'b1011101010;
    16'b0001000100010000: out_v[67] = 10'b0101101000;
    16'b0010000000010000: out_v[67] = 10'b0000110101;
    16'b0001000000000000: out_v[67] = 10'b1001001101;
    16'b0001000100000000: out_v[67] = 10'b0110011110;
    16'b0001000110010000: out_v[67] = 10'b1101010100;
    16'b0001000010000010: out_v[67] = 10'b0011110110;
    16'b0001000110010010: out_v[67] = 10'b1000001111;
    16'b0001000110010110: out_v[67] = 10'b1100011100;
    16'b0010010100010000: out_v[67] = 10'b1000011101;
    16'b0001000110000000: out_v[67] = 10'b0111011001;
    16'b0000000100000000: out_v[67] = 10'b1101000111;
    16'b0010000100000000: out_v[67] = 10'b1001010111;
    16'b0001000100010010: out_v[67] = 10'b0111001011;
    16'b0001000000000110: out_v[67] = 10'b1011001000;
    16'b0000010100010000: out_v[67] = 10'b1110001100;
    16'b0001000010000110: out_v[67] = 10'b0010011111;
    16'b0001010100010000: out_v[67] = 10'b0101111001;
    16'b0000000000010000: out_v[67] = 10'b0000100100;
    16'b0011000010000000: out_v[67] = 10'b0010101101;
    16'b0011000110010000: out_v[67] = 10'b1000011111;
    16'b0011000100000000: out_v[67] = 10'b0000001101;
    16'b0001000100010110: out_v[67] = 10'b0111011011;
    16'b0011000000010000: out_v[67] = 10'b1100000111;
    16'b0001000110000110: out_v[67] = 10'b0000010110;
    16'b0010000110010000: out_v[67] = 10'b1101011010;
    16'b0010000010000000: out_v[67] = 10'b1110000001;
    16'b0011010110010000: out_v[67] = 10'b1010101011;
    16'b0011110100010000: out_v[67] = 10'b0110011110;
    16'b0000010110010000: out_v[67] = 10'b0010100111;
    16'b0011010000000000: out_v[67] = 10'b0000011111;
    16'b0011010100000000: out_v[67] = 10'b0111011001;
    16'b0011010100010000: out_v[67] = 10'b1101010100;
    16'b0001000000000010: out_v[67] = 10'b0110000010;
    16'b0010000110000000: out_v[67] = 10'b1100101010;
    16'b0010010110000000: out_v[67] = 10'b1101101010;
    16'b0001010110010000: out_v[67] = 10'b1000011001;
    16'b0001110100010000: out_v[67] = 10'b0101100010;
    16'b0010010110010000: out_v[67] = 10'b0011011001;
    16'b0011010010000000: out_v[67] = 10'b0010011111;
    16'b0001110000000010: out_v[67] = 10'b1101011000;
    16'b0011110010000000: out_v[67] = 10'b0000110110;
    16'b0011110000000000: out_v[67] = 10'b1000000101;
    16'b0001110000000000: out_v[67] = 10'b1000001011;
    16'b0011100000000000: out_v[67] = 10'b0111110011;
    16'b0000110000000000: out_v[67] = 10'b1111101100;
    16'b0001100000000000: out_v[67] = 10'b0010111111;
    16'b0010110000000000: out_v[67] = 10'b0001011100;
    16'b0001100010000000: out_v[67] = 10'b1101010011;
    16'b0001110000000110: out_v[67] = 10'b1101110001;
    16'b0010010000000110: out_v[67] = 10'b1010100110;
    16'b0011110000000110: out_v[67] = 10'b0011100100;
    16'b0010110000000110: out_v[67] = 10'b0000100010;
    16'b0010000000000110: out_v[67] = 10'b0011110000;
    16'b0011010000000110: out_v[67] = 10'b0010110001;
    16'b0010110100010000: out_v[67] = 10'b0100110110;
    16'b0001110100000000: out_v[67] = 10'b1000111100;
    16'b0001100100010000: out_v[67] = 10'b0111100110;
    16'b0000110000010000: out_v[67] = 10'b0101110111;
    16'b0001010100000000: out_v[67] = 10'b0110110010;
    16'b0000110100000000: out_v[67] = 10'b1011011111;
    16'b0001010110000000: out_v[67] = 10'b1001010110;
    16'b0000010110000000: out_v[67] = 10'b1011110101;
    16'b0001100110010000: out_v[67] = 10'b0111110010;
    16'b0000010100000000: out_v[67] = 10'b0110010010;
    16'b0000100100010000: out_v[67] = 10'b1000111011;
    16'b0011000010000110: out_v[67] = 10'b1000110111;
    16'b0011110000000010: out_v[67] = 10'b0111001011;
    16'b0011110010000010: out_v[67] = 10'b1100111010;
    16'b0011000010000010: out_v[67] = 10'b0110110100;
    16'b0000010000000110: out_v[67] = 10'b1101001111;
    16'b0000010000000010: out_v[67] = 10'b1101100110;
    16'b0001110100010110: out_v[67] = 10'b1111011000;
    16'b0001010000000110: out_v[67] = 10'b1101111010;
    16'b0000000000000010: out_v[67] = 10'b0101011011;
    16'b0000110000000010: out_v[67] = 10'b1111100110;
    16'b0001110100010010: out_v[67] = 10'b1110110011;
    16'b0011000110110000: out_v[67] = 10'b1011011000;
    default: out_v[67] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000001101000: out_v[68] = 10'b1001010001;
    16'b0000000001101100: out_v[68] = 10'b1001011001;
    16'b0000000001001000: out_v[68] = 10'b0010100111;
    16'b0000000000101000: out_v[68] = 10'b0100110011;
    16'b0000000000000000: out_v[68] = 10'b1111100001;
    16'b0000000000001100: out_v[68] = 10'b0110100101;
    16'b0000000000001000: out_v[68] = 10'b0010100110;
    16'b0000000001001100: out_v[68] = 10'b0010100010;
    16'b0000000101101000: out_v[68] = 10'b0100110001;
    16'b0000010001101000: out_v[68] = 10'b0111000001;
    16'b0000000001000000: out_v[68] = 10'b1100101001;
    16'b0000010001000000: out_v[68] = 10'b0100000111;
    16'b0000000000101100: out_v[68] = 10'b0000111001;
    16'b0000000000100000: out_v[68] = 10'b1100110101;
    16'b0000000001000100: out_v[68] = 10'b1011100001;
    16'b0000010001100000: out_v[68] = 10'b0011010111;
    16'b0000010001001000: out_v[68] = 10'b1010101100;
    16'b0000000000000100: out_v[68] = 10'b1001001100;
    16'b0000010001000100: out_v[68] = 10'b0010001111;
    16'b0000010000100000: out_v[68] = 10'b1100010000;
    16'b0000000001100000: out_v[68] = 10'b1101110010;
    16'b0000010000000000: out_v[68] = 10'b1111000110;
    16'b0000000100000000: out_v[68] = 10'b0111001010;
    16'b0000000101000000: out_v[68] = 10'b0001101011;
    16'b0000000100100000: out_v[68] = 10'b0010000101;
    16'b0000000100100100: out_v[68] = 10'b0111000110;
    16'b0000000100000100: out_v[68] = 10'b0000101110;
    16'b0000000101001000: out_v[68] = 10'b1100110000;
    16'b1000000100000001: out_v[68] = 10'b1010110110;
    16'b0000010100000000: out_v[68] = 10'b1001001100;
    16'b0000010101000000: out_v[68] = 10'b0010011000;
    16'b1000010100100001: out_v[68] = 10'b0101010110;
    16'b0000000100001000: out_v[68] = 10'b1001010100;
    16'b0000010100100001: out_v[68] = 10'b0111000010;
    16'b0000000000100100: out_v[68] = 10'b0010111010;
    16'b0000010101100000: out_v[68] = 10'b0011101000;
    16'b0000010100000001: out_v[68] = 10'b1111110111;
    16'b1000000100100001: out_v[68] = 10'b1001000100;
    16'b0000010100100000: out_v[68] = 10'b1101000100;
    16'b1000010100000001: out_v[68] = 10'b1000110100;
    16'b0000000101100000: out_v[68] = 10'b0000011110;
    16'b0000000100100001: out_v[68] = 10'b1010110110;
    16'b0000000100101000: out_v[68] = 10'b0011100110;
    16'b1000010101100001: out_v[68] = 10'b1100010110;
    16'b0000010101001000: out_v[68] = 10'b0100011000;
    16'b0000010101101000: out_v[68] = 10'b0110100010;
    16'b0000010100001000: out_v[68] = 10'b0110110001;
    16'b0000010101000001: out_v[68] = 10'b0111101001;
    16'b1000010001001001: out_v[68] = 10'b1010110111;
    16'b1000000001001001: out_v[68] = 10'b0001011111;
    16'b0000010000001000: out_v[68] = 10'b0000111110;
    16'b0000010101000100: out_v[68] = 10'b0000111011;
    16'b0000000101000100: out_v[68] = 10'b1101001101;
    16'b1000000101001001: out_v[68] = 10'b1011001001;
    16'b1000010101001001: out_v[68] = 10'b0011101010;
    16'b1000010101000001: out_v[68] = 10'b1100111011;
    16'b0000010001001001: out_v[68] = 10'b0111100010;
    16'b0000010100101000: out_v[68] = 10'b1010111111;
    16'b0000000101001100: out_v[68] = 10'b1000100011;
    16'b0000000100001100: out_v[68] = 10'b1000011101;
    16'b0000010101100100: out_v[68] = 10'b0110010100;
    16'b0000000100101100: out_v[68] = 10'b1100110010;
    16'b0000000101101100: out_v[68] = 10'b1111110000;
    16'b0000010101001100: out_v[68] = 10'b1101101001;
    16'b0000010001001100: out_v[68] = 10'b1110110011;
    16'b0000010000101000: out_v[68] = 10'b0110101111;
    16'b0000000101100100: out_v[68] = 10'b0101100110;
    16'b0000010101101100: out_v[68] = 10'b0111110110;
    default: out_v[68] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100101100000000: out_v[69] = 10'b0100110101;
    16'b0100111101000000: out_v[69] = 10'b0101101011;
    16'b0100101001000000: out_v[69] = 10'b1010101001;
    16'b0100001100000000: out_v[69] = 10'b1001011000;
    16'b0100110101000000: out_v[69] = 10'b1110001011;
    16'b0100011100000100: out_v[69] = 10'b0001011110;
    16'b0100111100000000: out_v[69] = 10'b0100010111;
    16'b0100100100000000: out_v[69] = 10'b1110100001;
    16'b0100011100000000: out_v[69] = 10'b1111001101;
    16'b0000101100000000: out_v[69] = 10'b0101010011;
    16'b0000111100000000: out_v[69] = 10'b0010110010;
    16'b0100101100000100: out_v[69] = 10'b0111110101;
    16'b0100111001000000: out_v[69] = 10'b0110000111;
    16'b0100111101000100: out_v[69] = 10'b1011000101;
    16'b0100101101000000: out_v[69] = 10'b0000111010;
    16'b1100111100000000: out_v[69] = 10'b1011100111;
    16'b0100100101000000: out_v[69] = 10'b0100101010;
    16'b0100111100000100: out_v[69] = 10'b1011111010;
    16'b0000111001000000: out_v[69] = 10'b1111010100;
    16'b0100111100100000: out_v[69] = 10'b0011000011;
    16'b1100111100100000: out_v[69] = 10'b0100110011;
    16'b0100110001000000: out_v[69] = 10'b1110000010;
    16'b0100101000000000: out_v[69] = 10'b1010101110;
    16'b0000111101000000: out_v[69] = 10'b1000010011;
    16'b0100100001000000: out_v[69] = 10'b1001101111;
    16'b0100110100000000: out_v[69] = 10'b1100100001;
    16'b0000101001000000: out_v[69] = 10'b0000100111;
    16'b0100101101000100: out_v[69] = 10'b1111000000;
    16'b0100100100000100: out_v[69] = 10'b1001001111;
    16'b0100001001000000: out_v[69] = 10'b1101001011;
    16'b0100000100000000: out_v[69] = 10'b1111001000;
    16'b0100000000000100: out_v[69] = 10'b0000110011;
    16'b0000100100000100: out_v[69] = 10'b0011011010;
    16'b0000100100000000: out_v[69] = 10'b0010010110;
    16'b0000100000000100: out_v[69] = 10'b1000011011;
    16'b0000100101000100: out_v[69] = 10'b1100000011;
    16'b0100100000000100: out_v[69] = 10'b1111100100;
    16'b0000000100000000: out_v[69] = 10'b1100100000;
    16'b0100000100000100: out_v[69] = 10'b1100000001;
    16'b0100000000000000: out_v[69] = 10'b0010010011;
    16'b0100000000100100: out_v[69] = 10'b1101111000;
    16'b0000000000000000: out_v[69] = 10'b1001110111;
    16'b0000000000000100: out_v[69] = 10'b0011100111;
    16'b0000000000100100: out_v[69] = 10'b0101101110;
    16'b0000000000100000: out_v[69] = 10'b1001011010;
    16'b0000000100000100: out_v[69] = 10'b1110011100;
    16'b0100100001000101: out_v[69] = 10'b1110110011;
    16'b0000100001000100: out_v[69] = 10'b0111001100;
    16'b0100100001000100: out_v[69] = 10'b1010000000;
    16'b0100100000000101: out_v[69] = 10'b1111100110;
    16'b0100111000000100: out_v[69] = 10'b1100110100;
    16'b0100111001000101: out_v[69] = 10'b1111110110;
    16'b0100100000000001: out_v[69] = 10'b1000111110;
    16'b0100110100000100: out_v[69] = 10'b1011101100;
    16'b0100111001000100: out_v[69] = 10'b1000001100;
    16'b0100100101000101: out_v[69] = 10'b0001111110;
    16'b0100110000000100: out_v[69] = 10'b0011001111;
    16'b0100110001000100: out_v[69] = 10'b0100100111;
    16'b0100101001000101: out_v[69] = 10'b1011010111;
    16'b0100100101000100: out_v[69] = 10'b1110000100;
    16'b0100101001000100: out_v[69] = 10'b1110000101;
    16'b0000110000000100: out_v[69] = 10'b1001101111;
    16'b0100100001100100: out_v[69] = 10'b1001110101;
    16'b1100110000000100: out_v[69] = 10'b0111011011;
    16'b0000100000000101: out_v[69] = 10'b1101010011;
    16'b0100100001000001: out_v[69] = 10'b0011011011;
    16'b1100110100000100: out_v[69] = 10'b1111000011;
    16'b0000001101000100: out_v[69] = 10'b1000000101;
    16'b0100100000000000: out_v[69] = 10'b1001001001;
    16'b0100010000000100: out_v[69] = 10'b0001100100;
    16'b0000100101000101: out_v[69] = 10'b0110110101;
    16'b1000110000000100: out_v[69] = 10'b1110111110;
    16'b0000001100000100: out_v[69] = 10'b1110100101;
    16'b0100101000000101: out_v[69] = 10'b1110100100;
    16'b0000000101000100: out_v[69] = 10'b0000101011;
    16'b0100110101000100: out_v[69] = 10'b0111100101;
    16'b0100000001000100: out_v[69] = 10'b0000011010;
    16'b0100101000000100: out_v[69] = 10'b1000101101;
    16'b0000101101000100: out_v[69] = 10'b0001011011;
    16'b0100000000000101: out_v[69] = 10'b0110111100;
    16'b0100101001100000: out_v[69] = 10'b1111110011;
    16'b0000101100000001: out_v[69] = 10'b0011011000;
    16'b0100101101000001: out_v[69] = 10'b0101001010;
    16'b0100101001000001: out_v[69] = 10'b1011100000;
    16'b0000100000000000: out_v[69] = 10'b1100010100;
    16'b0000100101000000: out_v[69] = 10'b1101001101;
    16'b0000101101000001: out_v[69] = 10'b1111011111;
    16'b0000001101000000: out_v[69] = 10'b1110100001;
    16'b1100101001100000: out_v[69] = 10'b0010101000;
    16'b0000100001000000: out_v[69] = 10'b1000100101;
    16'b0100101000000001: out_v[69] = 10'b1111101100;
    16'b0100101001100001: out_v[69] = 10'b1111101001;
    16'b1100101001100001: out_v[69] = 10'b1111111001;
    16'b1100100001100000: out_v[69] = 10'b0111111011;
    16'b0000101101000000: out_v[69] = 10'b1000011011;
    16'b0100100001100000: out_v[69] = 10'b1111010100;
    16'b1100101001000000: out_v[69] = 10'b0111011011;
    16'b1100101101100000: out_v[69] = 10'b1011100000;
    16'b0100101100000001: out_v[69] = 10'b0110011111;
    16'b0100101101100000: out_v[69] = 10'b0100011010;
    16'b0100100101000001: out_v[69] = 10'b1010011011;
    16'b0100001000000100: out_v[69] = 10'b1000011001;
    16'b0100000001000000: out_v[69] = 10'b0000011001;
    16'b0100001001000100: out_v[69] = 10'b0001111010;
    16'b0000101100000100: out_v[69] = 10'b0011010000;
    16'b0000000001000100: out_v[69] = 10'b0001011000;
    16'b0000000001000000: out_v[69] = 10'b0001110001;
    16'b0000001000000100: out_v[69] = 10'b0011100010;
    16'b0000001001000000: out_v[69] = 10'b0101010100;
    16'b0000001000000000: out_v[69] = 10'b0010010110;
    16'b0000001001000100: out_v[69] = 10'b0001001010;
    16'b0000011000000100: out_v[69] = 10'b0101010011;
    16'b0100011000000100: out_v[69] = 10'b0000010011;
    16'b0100001000000000: out_v[69] = 10'b0001111010;
    16'b0000010000000100: out_v[69] = 10'b1010101001;
    16'b0000011001000100: out_v[69] = 10'b0001100111;
    16'b0100001100000100: out_v[69] = 10'b1001011001;
    16'b0000011001000000: out_v[69] = 10'b1011011011;
    16'b0000010100000100: out_v[69] = 10'b1010100110;
    16'b0000111100000100: out_v[69] = 10'b1011010000;
    16'b0000011100000100: out_v[69] = 10'b1100101111;
    16'b0000010001000000: out_v[69] = 10'b1101010010;
    16'b0100010100000100: out_v[69] = 10'b1101111100;
    16'b0100001101000000: out_v[69] = 10'b0010100000;
    16'b0100000101000000: out_v[69] = 10'b0001111110;
    16'b0100100100100000: out_v[69] = 10'b0101100110;
    16'b0100010100000000: out_v[69] = 10'b1100001110;
    16'b0000001001000101: out_v[69] = 10'b1011011001;
    16'b0000111101000100: out_v[69] = 10'b1001111011;
    16'b0000101000000100: out_v[69] = 10'b0100111100;
    16'b0000111001000100: out_v[69] = 10'b1011010110;
    16'b0000001000000101: out_v[69] = 10'b0111000010;
    16'b0000101001000100: out_v[69] = 10'b1100101011;
    16'b0000000000000101: out_v[69] = 10'b1101101011;
    16'b0000101000000000: out_v[69] = 10'b1001111010;
    16'b0000001100000000: out_v[69] = 10'b1010001100;
    16'b0100000101000100: out_v[69] = 10'b0110110011;
    16'b0000000101000000: out_v[69] = 10'b0111000000;
    16'b0100001101000100: out_v[69] = 10'b0110100011;
    16'b0100100100100100: out_v[69] = 10'b1001101111;
    16'b0100000100100100: out_v[69] = 10'b1101001100;
    default: out_v[69] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1001000010000001: out_v[70] = 10'b0000100101;
    16'b0001000010000001: out_v[70] = 10'b0000011101;
    16'b1011000110000001: out_v[70] = 10'b1111001101;
    16'b0001000000000001: out_v[70] = 10'b1101001000;
    16'b1001000010000000: out_v[70] = 10'b1100000111;
    16'b0000000000000000: out_v[70] = 10'b1011011001;
    16'b0001000010000000: out_v[70] = 10'b0010101001;
    16'b0001000110000001: out_v[70] = 10'b0010110011;
    16'b0001000000000000: out_v[70] = 10'b1111100011;
    16'b0011000000000001: out_v[70] = 10'b0011011011;
    16'b1001000110000001: out_v[70] = 10'b1000100100;
    16'b0000000010000001: out_v[70] = 10'b1001111100;
    16'b1011000010000001: out_v[70] = 10'b0110110011;
    16'b1000000010000000: out_v[70] = 10'b1011101010;
    16'b0000000000000001: out_v[70] = 10'b0000101110;
    16'b0000000010000000: out_v[70] = 10'b1110100001;
    16'b0011000010000001: out_v[70] = 10'b0110100011;
    16'b1000000010000001: out_v[70] = 10'b1001001000;
    16'b1001000010001001: out_v[70] = 10'b1001101111;
    16'b0000000100000001: out_v[70] = 10'b0101001011;
    16'b0011000110000001: out_v[70] = 10'b1010001101;
    16'b0001000010001001: out_v[70] = 10'b1011000111;
    16'b1000000000000001: out_v[70] = 10'b1100111001;
    16'b0011000100000001: out_v[70] = 10'b1111001110;
    16'b1011000010000000: out_v[70] = 10'b1001111000;
    16'b1000000000000000: out_v[70] = 10'b0111001011;
    16'b0000000000001001: out_v[70] = 10'b0000000110;
    16'b0000000000001000: out_v[70] = 10'b1011011011;
    16'b0000000010001000: out_v[70] = 10'b1111000010;
    16'b0001000000001000: out_v[70] = 10'b1100010100;
    16'b0001000010001000: out_v[70] = 10'b1111000000;
    16'b1001000000001000: out_v[70] = 10'b0001011110;
    16'b0000000000101000: out_v[70] = 10'b1010111001;
    16'b1001000010001000: out_v[70] = 10'b0101000100;
    16'b1000000000001000: out_v[70] = 10'b0100100011;
    16'b1001000110001000: out_v[70] = 10'b1110111100;
    16'b0010000000001001: out_v[70] = 10'b0101100111;
    16'b1000000010001000: out_v[70] = 10'b0101000110;
    16'b0000000100001001: out_v[70] = 10'b0110011011;
    16'b0001000000001001: out_v[70] = 10'b0010011001;
    16'b1011000000001000: out_v[70] = 10'b1111101111;
    16'b1011000100001000: out_v[70] = 10'b0010110111;
    16'b1001000000001001: out_v[70] = 10'b0010010010;
    16'b1001000100001000: out_v[70] = 10'b0010100111;
    16'b0000000100001000: out_v[70] = 10'b0111001100;
    16'b0010000100001001: out_v[70] = 10'b1001110111;
    16'b0001000100001000: out_v[70] = 10'b1101000111;
    16'b0010000000001000: out_v[70] = 10'b0011101111;
    16'b1000000100001000: out_v[70] = 10'b1001101111;
    16'b1001000000000000: out_v[70] = 10'b0000110110;
    16'b0001000110000000: out_v[70] = 10'b1011011001;
    16'b1001000110000000: out_v[70] = 10'b1110011010;
    16'b0000000100000000: out_v[70] = 10'b0111111001;
    16'b1001000000000001: out_v[70] = 10'b1001101000;
    16'b0000000110000000: out_v[70] = 10'b1011011111;
    16'b0000000010001001: out_v[70] = 10'b0010010010;
    16'b1000000000001001: out_v[70] = 10'b1100011010;
    16'b0001000010100000: out_v[70] = 10'b1011110110;
    16'b1001000010100001: out_v[70] = 10'b1110101011;
    16'b0000000110001000: out_v[70] = 10'b0011111110;
    16'b1000000010001001: out_v[70] = 10'b1101000010;
    default: out_v[70] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000000000001: out_v[71] = 10'b0001001110;
    16'b1100000000010000: out_v[71] = 10'b0001011011;
    16'b1100100000110001: out_v[71] = 10'b0001100011;
    16'b1100101000110001: out_v[71] = 10'b1100111001;
    16'b0000000000010001: out_v[71] = 10'b0111001010;
    16'b0000010000000000: out_v[71] = 10'b1010101101;
    16'b0100100000110001: out_v[71] = 10'b0110001100;
    16'b1100100000110000: out_v[71] = 10'b0010011111;
    16'b0100100000010000: out_v[71] = 10'b0010111111;
    16'b1100000000000000: out_v[71] = 10'b1011010011;
    16'b0100100000110000: out_v[71] = 10'b1110010001;
    16'b1100000000110001: out_v[71] = 10'b1111011010;
    16'b0000100000110001: out_v[71] = 10'b1110010011;
    16'b0000000000000000: out_v[71] = 10'b1101011100;
    16'b0101100000110000: out_v[71] = 10'b1110011011;
    16'b0100000000110001: out_v[71] = 10'b1111100110;
    16'b1100100000010001: out_v[71] = 10'b1011110111;
    16'b1000000000000000: out_v[71] = 10'b0010011001;
    16'b1001010000000000: out_v[71] = 10'b1111100011;
    16'b0000100000010001: out_v[71] = 10'b1010110010;
    16'b0100100000010001: out_v[71] = 10'b0110100111;
    16'b0000000000110001: out_v[71] = 10'b1110111111;
    16'b1100100000010000: out_v[71] = 10'b1111011111;
    16'b1100001000000000: out_v[71] = 10'b1101011011;
    16'b0101100000110001: out_v[71] = 10'b0011111000;
    16'b0100000000010001: out_v[71] = 10'b1111011110;
    16'b1100001000010000: out_v[71] = 10'b1101101110;
    16'b0101100000010000: out_v[71] = 10'b0101001111;
    16'b0101000000010000: out_v[71] = 10'b0001110001;
    16'b0100100000100001: out_v[71] = 10'b0110110001;
    16'b1100000000110000: out_v[71] = 10'b1101111010;
    16'b1000000000010000: out_v[71] = 10'b0101110011;
    16'b0100000000000000: out_v[71] = 10'b0110010101;
    16'b1000010000000000: out_v[71] = 10'b1100100001;
    16'b1100000000010001: out_v[71] = 10'b0010111110;
    16'b0000010000000001: out_v[71] = 10'b0000111111;
    16'b1100101000010000: out_v[71] = 10'b1111011100;
    16'b0100000000100001: out_v[71] = 10'b0010111011;
    16'b0001010000000000: out_v[71] = 10'b0011011110;
    16'b0000010000010001: out_v[71] = 10'b1010110111;
    16'b1000000000010001: out_v[71] = 10'b1001110001;
    16'b1100000000100001: out_v[71] = 10'b0010110101;
    16'b0100000000010000: out_v[71] = 10'b1111101011;
    16'b0000000000010000: out_v[71] = 10'b1100101010;
    16'b0001000000000000: out_v[71] = 10'b0011010111;
    16'b1001000000000000: out_v[71] = 10'b0100111111;
    16'b0001000000000001: out_v[71] = 10'b1011110100;
    16'b0001010000000001: out_v[71] = 10'b0011001100;
    16'b0000010000100000: out_v[71] = 10'b1000101100;
    16'b1001010000000001: out_v[71] = 10'b0011100100;
    16'b0001010000101000: out_v[71] = 10'b1111011110;
    16'b0001010000001000: out_v[71] = 10'b0001001100;
    16'b1000000000000001: out_v[71] = 10'b1111010111;
    16'b0001000000100001: out_v[71] = 10'b0001101100;
    16'b0101011000000000: out_v[71] = 10'b0111111100;
    16'b0001010000100000: out_v[71] = 10'b0100111101;
    16'b1001010000100000: out_v[71] = 10'b1001010111;
    16'b0001010000001001: out_v[71] = 10'b1011011101;
    16'b1001010000100001: out_v[71] = 10'b1010010111;
    16'b0001000000001001: out_v[71] = 10'b1111111111;
    16'b0001010000100001: out_v[71] = 10'b1011001011;
    16'b0001000000100000: out_v[71] = 10'b1000000101;
    16'b0001011000001000: out_v[71] = 10'b1000111011;
    16'b0000000000100000: out_v[71] = 10'b0111110110;
    16'b1001000000000001: out_v[71] = 10'b1000110110;
    16'b0001000000101000: out_v[71] = 10'b1011000011;
    16'b1000010000000001: out_v[71] = 10'b0001011010;
    16'b0000000000100001: out_v[71] = 10'b0101101110;
    16'b0001011000100000: out_v[71] = 10'b1111010111;
    16'b0001000000101001: out_v[71] = 10'b0100001110;
    16'b0001011000000001: out_v[71] = 10'b0111100111;
    16'b0001011000101000: out_v[71] = 10'b0111110011;
    16'b1000010000100000: out_v[71] = 10'b1001001111;
    16'b0001011000001001: out_v[71] = 10'b0110010111;
    16'b0000000000001001: out_v[71] = 10'b1010100111;
    16'b0000010000001000: out_v[71] = 10'b1101100000;
    16'b0001010000101001: out_v[71] = 10'b0111100101;
    16'b0001011000000000: out_v[71] = 10'b0001001111;
    16'b1000001000000000: out_v[71] = 10'b1101011110;
    16'b1000011000100001: out_v[71] = 10'b1011111000;
    16'b0000010000100001: out_v[71] = 10'b1000101010;
    16'b1000010000110001: out_v[71] = 10'b1011111011;
    16'b1000010000100001: out_v[71] = 10'b1010011011;
    16'b1000011000000000: out_v[71] = 10'b0100100010;
    16'b1000011000000001: out_v[71] = 10'b1110000010;
    16'b0000011000000000: out_v[71] = 10'b1011110110;
    16'b1000010000010000: out_v[71] = 10'b0110001011;
    16'b0000010000110001: out_v[71] = 10'b0010111011;
    16'b1000010000010001: out_v[71] = 10'b1101100111;
    16'b1000000000100001: out_v[71] = 10'b1001001001;
    16'b0000110000110001: out_v[71] = 10'b0010110001;
    16'b1000110000110001: out_v[71] = 10'b0110100010;
    16'b0001010000010001: out_v[71] = 10'b1100000011;
    16'b0001110000010001: out_v[71] = 10'b0101010001;
    16'b0000010000010000: out_v[71] = 10'b1000101011;
    16'b0000110000010001: out_v[71] = 10'b0110010110;
    16'b0001010000010000: out_v[71] = 10'b1100100111;
    16'b0001110000010000: out_v[71] = 10'b1010111101;
    16'b1001110000010000: out_v[71] = 10'b0011110100;
    16'b0000110000010000: out_v[71] = 10'b1101010010;
    16'b0101010000010000: out_v[71] = 10'b1101101010;
    16'b0100110000010000: out_v[71] = 10'b1101010011;
    16'b0000110000110000: out_v[71] = 10'b0100110011;
    16'b0101110000010000: out_v[71] = 10'b0010011000;
    16'b0100110000010001: out_v[71] = 10'b0001111110;
    16'b0001110000110000: out_v[71] = 10'b0111010010;
    16'b1001010000010000: out_v[71] = 10'b0111011101;
    16'b0000110000000001: out_v[71] = 10'b0000011011;
    16'b0001000000010000: out_v[71] = 10'b0111010000;
    16'b1001000000010000: out_v[71] = 10'b0011111110;
    16'b1000110000010001: out_v[71] = 10'b1011111000;
    16'b1000100000010001: out_v[71] = 10'b1011110110;
    16'b1000100000010000: out_v[71] = 10'b0101100011;
    16'b0001100000010001: out_v[71] = 10'b0101101010;
    16'b0000100000010000: out_v[71] = 10'b0010101001;
    16'b1000110000010000: out_v[71] = 10'b1011101010;
    16'b0001010000111001: out_v[71] = 10'b1011010101;
    16'b0101110000110001: out_v[71] = 10'b1010101011;
    16'b0001010000110000: out_v[71] = 10'b1111100000;
    16'b0001000000001000: out_v[71] = 10'b1001010100;
    16'b0000110000111001: out_v[71] = 10'b0011011110;
    16'b0001010000111000: out_v[71] = 10'b1000110111;
    16'b0101110000111000: out_v[71] = 10'b1000110111;
    16'b0101110000110000: out_v[71] = 10'b0111010011;
    16'b0101010000000000: out_v[71] = 10'b0110111110;
    16'b0001110000111001: out_v[71] = 10'b0011111011;
    16'b0000010000001001: out_v[71] = 10'b0010110010;
    16'b0001010000011000: out_v[71] = 10'b1111001011;
    16'b0101010000001000: out_v[71] = 10'b1000101110;
    16'b0001110000110001: out_v[71] = 10'b1110001010;
    16'b0101010000011000: out_v[71] = 10'b0011101001;
    16'b0000010000101001: out_v[71] = 10'b1100100010;
    16'b0001010000110001: out_v[71] = 10'b0111001111;
    16'b0000000000001000: out_v[71] = 10'b1100111001;
    16'b0101110000111001: out_v[71] = 10'b1101010010;
    16'b0000010000111001: out_v[71] = 10'b1011000100;
    16'b0101010000111000: out_v[71] = 10'b0110111010;
    16'b0101010000110001: out_v[71] = 10'b1000111011;
    16'b0101010000110000: out_v[71] = 10'b1111101010;
    16'b1101110000010000: out_v[71] = 10'b0010010010;
    16'b1001010100000000: out_v[71] = 10'b1111000011;
    16'b0000110000000000: out_v[71] = 10'b1100100111;
    16'b1101010000000000: out_v[71] = 10'b1100010011;
    16'b0100010000000000: out_v[71] = 10'b0110100100;
    16'b1101010100000000: out_v[71] = 10'b1010100010;
    16'b1100010000000000: out_v[71] = 10'b0101011100;
    16'b0001000000010001: out_v[71] = 10'b0110100110;
    16'b1101010000010000: out_v[71] = 10'b1101011011;
    16'b1001010000010001: out_v[71] = 10'b0001011110;
    16'b0001110000000001: out_v[71] = 10'b0001101111;
    default: out_v[71] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000000001000: out_v[72] = 10'b1000101101;
    16'b0100001000010010: out_v[72] = 10'b1110111111;
    16'b0100001000010101: out_v[72] = 10'b1100000011;
    16'b0000001000001100: out_v[72] = 10'b1110111110;
    16'b0010001000011100: out_v[72] = 10'b0000000111;
    16'b0100001000010001: out_v[72] = 10'b1111010011;
    16'b0010001000010010: out_v[72] = 10'b1111001001;
    16'b0100000000010000: out_v[72] = 10'b1100011011;
    16'b0100001000010100: out_v[72] = 10'b1100011111;
    16'b0100001000000001: out_v[72] = 10'b0111110000;
    16'b0010001000011000: out_v[72] = 10'b1101010001;
    16'b0000001000011100: out_v[72] = 10'b1001010101;
    16'b0100001000010000: out_v[72] = 10'b0001111100;
    16'b0010001100011100: out_v[72] = 10'b1100111000;
    16'b0000001000011000: out_v[72] = 10'b1101101101;
    16'b0000001000010110: out_v[72] = 10'b1110111001;
    16'b0000000000000000: out_v[72] = 10'b0111001000;
    16'b0000001000000001: out_v[72] = 10'b0001111110;
    16'b0000001000010000: out_v[72] = 10'b0101101011;
    16'b0010001000010000: out_v[72] = 10'b0111010000;
    16'b0010001000010100: out_v[72] = 10'b0100100111;
    16'b0000001000011101: out_v[72] = 10'b1111011101;
    16'b0100001000010110: out_v[72] = 10'b1101110010;
    16'b0100000000000001: out_v[72] = 10'b1000001011;
    16'b0000001000010010: out_v[72] = 10'b1001101001;
    16'b0000001000010100: out_v[72] = 10'b1110101010;
    16'b0000001000000100: out_v[72] = 10'b1000110111;
    16'b0000001000001001: out_v[72] = 10'b0010110111;
    16'b0000001000001000: out_v[72] = 10'b0111110011;
    16'b0010001000010110: out_v[72] = 10'b1110001001;
    16'b0000000000000100: out_v[72] = 10'b1111010001;
    16'b0100001000000101: out_v[72] = 10'b1110101101;
    16'b0010001000011010: out_v[72] = 10'b0010111010;
    16'b0010000000001000: out_v[72] = 10'b1010000111;
    16'b0100000000000000: out_v[72] = 10'b1101011001;
    16'b0100001000011001: out_v[72] = 10'b1011101001;
    16'b0000000000000001: out_v[72] = 10'b1001001110;
    16'b0000000000001001: out_v[72] = 10'b0110110011;
    16'b0000000000001100: out_v[72] = 10'b1011100111;
    16'b0000001000000101: out_v[72] = 10'b1010110100;
    16'b0110001000010000: out_v[72] = 10'b0100110100;
    16'b0000001000011001: out_v[72] = 10'b1000011101;
    16'b0010001100011000: out_v[72] = 10'b0011011001;
    16'b0000001000000000: out_v[72] = 10'b0110101101;
    16'b0000000100001000: out_v[72] = 10'b1100110011;
    16'b0000000100010000: out_v[72] = 10'b0001111100;
    16'b0000001100010000: out_v[72] = 10'b0000010101;
    16'b0000000100000100: out_v[72] = 10'b1011011011;
    16'b0000001100010100: out_v[72] = 10'b0110110011;
    16'b0000000100000000: out_v[72] = 10'b1000000011;
    16'b0000001100000000: out_v[72] = 10'b1110001110;
    16'b0000001100000100: out_v[72] = 10'b1011100111;
    16'b0000000100001100: out_v[72] = 10'b0001111010;
    16'b0010000100010000: out_v[72] = 10'b1000100110;
    16'b0000001100011000: out_v[72] = 10'b0111100000;
    16'b0010001100010100: out_v[72] = 10'b1110101000;
    16'b0000000100001010: out_v[72] = 10'b1011001011;
    16'b0000001100011100: out_v[72] = 10'b1001011110;
    16'b0000001100001100: out_v[72] = 10'b1100111010;
    16'b0000000000010000: out_v[72] = 10'b0001111110;
    16'b0010001100010000: out_v[72] = 10'b1000001011;
    16'b0000001100011001: out_v[72] = 10'b1001000111;
    16'b0000001100010001: out_v[72] = 10'b1001100101;
    16'b0010001100010001: out_v[72] = 10'b0001011111;
    16'b0000001100010101: out_v[72] = 10'b1011101011;
    16'b0010000000001100: out_v[72] = 10'b1000100010;
    16'b0010000000001101: out_v[72] = 10'b0101010011;
    16'b0000001100011101: out_v[72] = 10'b0000100110;
    16'b0010001000011101: out_v[72] = 10'b1011000110;
    16'b0110000100001000: out_v[72] = 10'b0011101111;
    16'b0010000000000000: out_v[72] = 10'b1011100000;
    16'b0010000000011000: out_v[72] = 10'b1000001010;
    16'b0010001000010101: out_v[72] = 10'b1000100011;
    16'b0010001000011001: out_v[72] = 10'b0110100010;
    16'b0010000000011101: out_v[72] = 10'b0100101011;
    16'b0010000000001001: out_v[72] = 10'b0010110000;
    16'b0010000100001000: out_v[72] = 10'b1010000101;
    16'b0010001000010001: out_v[72] = 10'b0100010100;
    16'b0010001100011001: out_v[72] = 10'b0110101111;
    16'b0010000000011001: out_v[72] = 10'b1001101110;
    16'b0000000100011101: out_v[72] = 10'b1001111011;
    16'b0010000000011100: out_v[72] = 10'b0011010010;
    16'b0000001000010101: out_v[72] = 10'b1111011101;
    16'b0010001100011101: out_v[72] = 10'b1111111001;
    16'b0110000000001000: out_v[72] = 10'b0101000110;
    16'b0010000100011000: out_v[72] = 10'b0011111001;
    16'b0010000100001100: out_v[72] = 10'b0110011010;
    16'b0000000100011001: out_v[72] = 10'b0110111000;
    16'b0000000100011000: out_v[72] = 10'b1101110111;
    16'b0010000000000100: out_v[72] = 10'b0101111110;
    16'b0110001000011000: out_v[72] = 10'b1010111110;
    16'b0010001100000000: out_v[72] = 10'b1000000000;
    16'b0010000000000001: out_v[72] = 10'b0101111110;
    16'b1010001100010100: out_v[72] = 10'b1110101011;
    16'b1000001100010100: out_v[72] = 10'b1111011010;
    16'b0010000100000000: out_v[72] = 10'b1011010010;
    16'b0000000100000001: out_v[72] = 10'b0010011101;
    16'b1010001100010000: out_v[72] = 10'b0100011110;
    16'b1000001100010000: out_v[72] = 10'b1101001111;
    16'b1010001100011100: out_v[72] = 10'b1010011011;
    16'b0010000100000001: out_v[72] = 10'b1101011011;
    16'b0000000100001001: out_v[72] = 10'b1111110110;
    16'b0010001100001001: out_v[72] = 10'b0010011011;
    16'b0000001100000001: out_v[72] = 10'b0011110010;
    16'b0010001100001000: out_v[72] = 10'b0100110100;
    16'b0010001100000100: out_v[72] = 10'b1110110111;
    16'b0010000100001001: out_v[72] = 10'b0100011111;
    16'b0010001100000001: out_v[72] = 10'b1001001011;
    16'b1010001100011000: out_v[72] = 10'b0111001011;
    16'b0010000100000100: out_v[72] = 10'b1100100010;
    16'b0010001100010101: out_v[72] = 10'b1000111011;
    16'b0110001100011000: out_v[72] = 10'b1010010010;
    16'b0010000000001010: out_v[72] = 10'b1101110010;
    16'b0010000000010000: out_v[72] = 10'b0111110001;
    16'b0110000000011000: out_v[72] = 10'b0110111011;
    16'b0010000000011010: out_v[72] = 10'b0101100010;
    16'b0010001100011010: out_v[72] = 10'b0001111010;
    16'b0010001100010010: out_v[72] = 10'b0000110001;
    16'b0000000000011010: out_v[72] = 10'b0011111011;
    16'b0010000100010010: out_v[72] = 10'b0011101100;
    16'b0000001000011010: out_v[72] = 10'b0000101110;
    16'b0010000000000010: out_v[72] = 10'b1000010101;
    16'b0000000000010010: out_v[72] = 10'b1011101111;
    16'b0100000100000001: out_v[72] = 10'b0110110100;
    16'b0000000000001010: out_v[72] = 10'b0101110110;
    16'b0000001001011010: out_v[72] = 10'b1010111111;
    16'b0010000000000011: out_v[72] = 10'b1101110010;
    16'b0000001100010010: out_v[72] = 10'b0101110001;
    16'b0000000000011000: out_v[72] = 10'b0010100101;
    16'b0010001000111100: out_v[72] = 10'b1110101011;
    16'b0100001100010000: out_v[72] = 10'b1001011011;
    16'b0010001000001100: out_v[72] = 10'b1011000011;
    16'b0110001000111100: out_v[72] = 10'b1110110011;
    16'b0110001000011001: out_v[72] = 10'b1110100001;
    16'b0000001000111100: out_v[72] = 10'b1000111101;
    16'b0010001100111100: out_v[72] = 10'b1111001110;
    16'b0100001100011000: out_v[72] = 10'b1010011011;
    16'b0000001100111100: out_v[72] = 10'b1111001100;
    16'b0110001000011100: out_v[72] = 10'b1010011010;
    16'b0100001000011000: out_v[72] = 10'b0111001010;
    16'b0010001000111000: out_v[72] = 10'b0010011010;
    16'b0010001000110100: out_v[72] = 10'b0110011101;
    16'b0010000000111100: out_v[72] = 10'b1101100011;
    16'b0100001100011001: out_v[72] = 10'b0011001001;
    16'b0010001100001100: out_v[72] = 10'b1100000010;
    16'b0000001100011010: out_v[72] = 10'b0101011000;
    16'b0000001100001000: out_v[72] = 10'b0110011011;
    16'b0010001100001101: out_v[72] = 10'b1111010011;
    16'b0010000100001010: out_v[72] = 10'b0100011001;
    16'b0000000100011010: out_v[72] = 10'b0110000011;
    16'b0010100000001000: out_v[72] = 10'b1111100111;
    16'b0010100000001001: out_v[72] = 10'b1000100101;
    16'b0010100100001000: out_v[72] = 10'b1100101000;
    16'b0010100100001001: out_v[72] = 10'b1101000101;
    default: out_v[72] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010001000011000: out_v[73] = 10'b0110010111;
    16'b0010001000001000: out_v[73] = 10'b0001101100;
    16'b0010000000001000: out_v[73] = 10'b0010000011;
    16'b0110000000011000: out_v[73] = 10'b0010011101;
    16'b0010000000011000: out_v[73] = 10'b0010011111;
    16'b0000000000001000: out_v[73] = 10'b0010101010;
    16'b0000000000011000: out_v[73] = 10'b1111000011;
    16'b0100000000010000: out_v[73] = 10'b0001011111;
    16'b0110001000011000: out_v[73] = 10'b1110000011;
    16'b0110001000010000: out_v[73] = 10'b0111001010;
    16'b0000000000001001: out_v[73] = 10'b0110101000;
    16'b0110001000011001: out_v[73] = 10'b0010101111;
    16'b0010000000011001: out_v[73] = 10'b1011110010;
    16'b0010001000000000: out_v[73] = 10'b0011110101;
    16'b0010000000000000: out_v[73] = 10'b0011011000;
    16'b0010000000001001: out_v[73] = 10'b1111001100;
    16'b0110000000011001: out_v[73] = 10'b1101010010;
    16'b0010000000100001: out_v[73] = 10'b1101001011;
    16'b0010001000000001: out_v[73] = 10'b0011101001;
    16'b0110000000010000: out_v[73] = 10'b1101010111;
    16'b0000000000010000: out_v[73] = 10'b0000101111;
    16'b0010000000010000: out_v[73] = 10'b1101110011;
    16'b0110000000111001: out_v[73] = 10'b1111011011;
    16'b0010000000111001: out_v[73] = 10'b1100010011;
    16'b0100000000011000: out_v[73] = 10'b1001010100;
    16'b0010001000001001: out_v[73] = 10'b1000101001;
    16'b0010000000000001: out_v[73] = 10'b0110001110;
    16'b0010001000011001: out_v[73] = 10'b1101101110;
    16'b0100000000011001: out_v[73] = 10'b1000011011;
    16'b0010000000101001: out_v[73] = 10'b0001101100;
    16'b0100000000111001: out_v[73] = 10'b0110110011;
    16'b0100001000011000: out_v[73] = 10'b0010111011;
    16'b0000000000011001: out_v[73] = 10'b1101000000;
    16'b0100000000000000: out_v[73] = 10'b1001101110;
    16'b0000000000000000: out_v[73] = 10'b0010111000;
    16'b0000001000000000: out_v[73] = 10'b1111110000;
    16'b0110000000000000: out_v[73] = 10'b0110101100;
    16'b0100001000000000: out_v[73] = 10'b0111011001;
    16'b0000000000000001: out_v[73] = 10'b0000000011;
    16'b0000000000100000: out_v[73] = 10'b1100111000;
    16'b0100000000100001: out_v[73] = 10'b0000011011;
    16'b0100000000110001: out_v[73] = 10'b1001010100;
    16'b0100000000111000: out_v[73] = 10'b1010110110;
    16'b0000000000100001: out_v[73] = 10'b0100101100;
    16'b0110000000110001: out_v[73] = 10'b1110000111;
    16'b0010000000100000: out_v[73] = 10'b1010101011;
    16'b0010000000101000: out_v[73] = 10'b0010101111;
    16'b0100000000010001: out_v[73] = 10'b0011101001;
    16'b0110000000010001: out_v[73] = 10'b0010000111;
    16'b0100000000110000: out_v[73] = 10'b0000111110;
    16'b0110000000111000: out_v[73] = 10'b1011000101;
    16'b0100000000100000: out_v[73] = 10'b0110110111;
    16'b0110000000110000: out_v[73] = 10'b0011010100;
    16'b0000000000101000: out_v[73] = 10'b1101001100;
    16'b0100000000101000: out_v[73] = 10'b1001100111;
    16'b0100000000001000: out_v[73] = 10'b1100010011;
    16'b0100000000000001: out_v[73] = 10'b0010001110;
    16'b0000001000001000: out_v[73] = 10'b1010100110;
    16'b0000001000101000: out_v[73] = 10'b1011101110;
    16'b0000001000100001: out_v[73] = 10'b0001110110;
    16'b0000001000001001: out_v[73] = 10'b0001011111;
    16'b0000001000101001: out_v[73] = 10'b1011110110;
    16'b0000000000101001: out_v[73] = 10'b0001101001;
    16'b0000001000100000: out_v[73] = 10'b0011010111;
    16'b0000001000000001: out_v[73] = 10'b1010101111;
    16'b0010001000101000: out_v[73] = 10'b0111100101;
    16'b0010001000101001: out_v[73] = 10'b0001101010;
    16'b0010001000100000: out_v[73] = 10'b1101111010;
    16'b0000000000000010: out_v[73] = 10'b0000011101;
    16'b0100001000010000: out_v[73] = 10'b1110001000;
    16'b0001000000000000: out_v[73] = 10'b1011110010;
    16'b0010000000000010: out_v[73] = 10'b1010000101;
    16'b0010000000001010: out_v[73] = 10'b1000100011;
    16'b0110000000010010: out_v[73] = 10'b0110001011;
    16'b0010001000000010: out_v[73] = 10'b0111101100;
    16'b0110001000010010: out_v[73] = 10'b0101100011;
    16'b0010000000010010: out_v[73] = 10'b0100111111;
    16'b0100000000001001: out_v[73] = 10'b1111011011;
    16'b0100010000011000: out_v[73] = 10'b1010110100;
    16'b0100010000010000: out_v[73] = 10'b1111100110;
    16'b0000000000111000: out_v[73] = 10'b1010110110;
    16'b0000010000001000: out_v[73] = 10'b0111100010;
    16'b0000010000011000: out_v[73] = 10'b1001000111;
    16'b0100010000001000: out_v[73] = 10'b1111110011;
    16'b0100010000000000: out_v[73] = 10'b0111001100;
    16'b0100010000011001: out_v[73] = 10'b1101110111;
    16'b0010001001000000: out_v[73] = 10'b0001001010;
    16'b0000000100000000: out_v[73] = 10'b1000111001;
    16'b0110001000010001: out_v[73] = 10'b0101010010;
    16'b0110001000000000: out_v[73] = 10'b0001011111;
    16'b0100001000010010: out_v[73] = 10'b0101011111;
    16'b0100000000010010: out_v[73] = 10'b1101001101;
    16'b0100001000011001: out_v[73] = 10'b0110100111;
    16'b0110000001011001: out_v[73] = 10'b1001000010;
    16'b0100000001011001: out_v[73] = 10'b1011001110;
    default: out_v[73] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000010000000000: out_v[74] = 10'b0010010101;
    16'b0010010000000000: out_v[74] = 10'b0010010101;
    16'b0010010001001000: out_v[74] = 10'b1001001011;
    16'b0010010001000000: out_v[74] = 10'b1000010101;
    16'b0000010001001000: out_v[74] = 10'b1011000101;
    16'b0010000000000000: out_v[74] = 10'b1001001100;
    16'b0000000001000000: out_v[74] = 10'b0000111101;
    16'b0000000000000000: out_v[74] = 10'b0011100111;
    16'b0010010100000000: out_v[74] = 10'b0011101010;
    16'b0000010110000000: out_v[74] = 10'b1100011001;
    16'b0010010000001000: out_v[74] = 10'b0010010101;
    16'b0010010101000000: out_v[74] = 10'b0100011001;
    16'b0000010001000000: out_v[74] = 10'b1001011100;
    16'b0000000001001000: out_v[74] = 10'b0011011011;
    16'b0010000001000000: out_v[74] = 10'b1001110001;
    16'b0000010100000000: out_v[74] = 10'b1101001010;
    16'b0000000100000000: out_v[74] = 10'b1011111110;
    16'b0010000001001000: out_v[74] = 10'b1101010011;
    16'b0000010010000000: out_v[74] = 10'b1100100100;
    16'b0000000010000000: out_v[74] = 10'b0001011010;
    16'b0010010101001000: out_v[74] = 10'b1010000111;
    16'b0000000110000000: out_v[74] = 10'b0110110010;
    16'b0000000101000000: out_v[74] = 10'b1000101110;
    16'b0000000111000000: out_v[74] = 10'b1101010001;
    16'b0010010010000000: out_v[74] = 10'b1000110100;
    16'b0000010000001000: out_v[74] = 10'b0000001100;
    16'b0000000011000000: out_v[74] = 10'b1000110101;
    16'b0000000111001000: out_v[74] = 10'b1101000000;
    16'b0010010110000000: out_v[74] = 10'b0011011011;
    16'b0000010011000000: out_v[74] = 10'b0111000110;
    16'b0000010111000000: out_v[74] = 10'b1101010100;
    16'b0010000110000000: out_v[74] = 10'b1000010110;
    16'b0000000101001000: out_v[74] = 10'b1000110010;
    16'b0000010101000000: out_v[74] = 10'b1011001101;
    16'b0010000010000000: out_v[74] = 10'b0010000111;
    16'b0010000100000000: out_v[74] = 10'b0010111000;
    16'b0010000111000000: out_v[74] = 10'b0011101010;
    16'b1010000101000000: out_v[74] = 10'b1100011010;
    16'b1010000111000000: out_v[74] = 10'b1011101001;
    16'b0010000101000000: out_v[74] = 10'b0000100100;
    16'b1000000101000000: out_v[74] = 10'b0001101100;
    16'b1000000111000000: out_v[74] = 10'b0000101011;
    16'b0010010111000000: out_v[74] = 10'b1100011000;
    16'b0010000101001000: out_v[74] = 10'b0010101001;
    16'b0010000111001000: out_v[74] = 10'b0101111011;
    16'b0000010010001000: out_v[74] = 10'b1100111011;
    16'b0000000110001000: out_v[74] = 10'b0101011001;
    16'b0000010011001000: out_v[74] = 10'b0101000000;
    16'b0000000010001000: out_v[74] = 10'b1100100111;
    16'b0010010011001000: out_v[74] = 10'b1010010010;
    16'b0100010010000000: out_v[74] = 10'b1101010100;
    16'b0100000100000000: out_v[74] = 10'b0010101010;
    16'b0100000010000000: out_v[74] = 10'b0100101010;
    16'b0000000011001000: out_v[74] = 10'b0101100010;
    16'b0010000011000000: out_v[74] = 10'b1001100100;
    16'b0000000010100000: out_v[74] = 10'b0110101011;
    16'b0000000110100000: out_v[74] = 10'b1011101101;
    16'b0010000001100000: out_v[74] = 10'b0111000101;
    16'b0010000000100000: out_v[74] = 10'b0101100010;
    16'b0000000000100000: out_v[74] = 10'b1111001111;
    16'b0010000110100000: out_v[74] = 10'b1100100111;
    16'b0010000010100000: out_v[74] = 10'b1111101001;
    16'b0010000011100000: out_v[74] = 10'b1110110011;
    16'b0010000111100000: out_v[74] = 10'b1110101010;
    16'b0000010100001000: out_v[74] = 10'b0110010110;
    16'b0000000000001000: out_v[74] = 10'b1001000100;
    16'b0000000100001000: out_v[74] = 10'b0111100000;
    16'b0000010111001000: out_v[74] = 10'b1101100110;
    16'b0010010111001000: out_v[74] = 10'b1011001010;
    16'b0000010110001000: out_v[74] = 10'b1001011100;
    default: out_v[74] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001010000000001: out_v[75] = 10'b1010010001;
    16'b0011010000000001: out_v[75] = 10'b0000100001;
    16'b0011000000000000: out_v[75] = 10'b1001000011;
    16'b0000010000000000: out_v[75] = 10'b0000000011;
    16'b0001000000000000: out_v[75] = 10'b0010011100;
    16'b0001010000000000: out_v[75] = 10'b0000000001;
    16'b0010010000000000: out_v[75] = 10'b1000000111;
    16'b0010010000000001: out_v[75] = 10'b0010110001;
    16'b0010000000000000: out_v[75] = 10'b0010110011;
    16'b0011110000000001: out_v[75] = 10'b1000010111;
    16'b0011010000000000: out_v[75] = 10'b1000100001;
    16'b0011000000000001: out_v[75] = 10'b0110000110;
    16'b0011110000000000: out_v[75] = 10'b0011100110;
    16'b0001010010000000: out_v[75] = 10'b0110001100;
    16'b0011110000000100: out_v[75] = 10'b1000111011;
    16'b0011010000010001: out_v[75] = 10'b0101000110;
    16'b0011010010000001: out_v[75] = 10'b1000001111;
    16'b0000000000000000: out_v[75] = 10'b0101001101;
    16'b0011010000000100: out_v[75] = 10'b0110011001;
    16'b0000010010000000: out_v[75] = 10'b1101101001;
    16'b0011010010010001: out_v[75] = 10'b1001011010;
    16'b0011000000010001: out_v[75] = 10'b1000000111;
    16'b0001010010010000: out_v[75] = 10'b0010011010;
    16'b0000000010010000: out_v[75] = 10'b0000001111;
    16'b0000010000010000: out_v[75] = 10'b1001101010;
    16'b0000000000010000: out_v[75] = 10'b0100010110;
    16'b0000000010000000: out_v[75] = 10'b1001001001;
    16'b0001000010000000: out_v[75] = 10'b0000111110;
    16'b0001000010010000: out_v[75] = 10'b1100101110;
    16'b0000010010010000: out_v[75] = 10'b0010000111;
    16'b0000110010010000: out_v[75] = 10'b1110110101;
    16'b0000110010010100: out_v[75] = 10'b1110110111;
    16'b0001100010010000: out_v[75] = 10'b1110101001;
    16'b0001110010000100: out_v[75] = 10'b0110010111;
    16'b0000110010000000: out_v[75] = 10'b0010100001;
    16'b0001110010010100: out_v[75] = 10'b1001110011;
    16'b0011000010010001: out_v[75] = 10'b1000110111;
    16'b0001110000000000: out_v[75] = 10'b0001011010;
    16'b0010000000010001: out_v[75] = 10'b0100011110;
    16'b0001000010010100: out_v[75] = 10'b0001000111;
    16'b0000100010010000: out_v[75] = 10'b0111100101;
    16'b0011110000010001: out_v[75] = 10'b1111010110;
    16'b0000110010000100: out_v[75] = 10'b1010111111;
    16'b0001100010010100: out_v[75] = 10'b1001100110;
    16'b0000000010010100: out_v[75] = 10'b0110010111;
    16'b0001110010010000: out_v[75] = 10'b1110111011;
    16'b0001110010000000: out_v[75] = 10'b0101100010;
    16'b0001010010010100: out_v[75] = 10'b1010000111;
    16'b0000110000000100: out_v[75] = 10'b0111000111;
    16'b0010000010010001: out_v[75] = 10'b0011011000;
    16'b0000100010010100: out_v[75] = 10'b1100000100;
    16'b0011000010010000: out_v[75] = 10'b1111010111;
    16'b0000110000000000: out_v[75] = 10'b0000111101;
    16'b0000100000010000: out_v[75] = 10'b1000100101;
    16'b0001010000010000: out_v[75] = 10'b0110111000;
    16'b0000100010000000: out_v[75] = 10'b0101011011;
    16'b0011010010000000: out_v[75] = 10'b0111001000;
    16'b0001010010000001: out_v[75] = 10'b1110001011;
    16'b0001110010000001: out_v[75] = 10'b1011110011;
    16'b0000010000000001: out_v[75] = 10'b0001110010;
    16'b0000110000000001: out_v[75] = 10'b0010110011;
    16'b0000110010000001: out_v[75] = 10'b1000110100;
    16'b0000110010000010: out_v[75] = 10'b1010111011;
    16'b0010010010010001: out_v[75] = 10'b0111010000;
    16'b0001010010010001: out_v[75] = 10'b0110111101;
    16'b0011010010010000: out_v[75] = 10'b1101010000;
    16'b0010000010000001: out_v[75] = 10'b1010001011;
    16'b0001000010010001: out_v[75] = 10'b0000010111;
    16'b0010010010000001: out_v[75] = 10'b1110001110;
    16'b0011000010000001: out_v[75] = 10'b1000011010;
    16'b0001000000010000: out_v[75] = 10'b1101111000;
    16'b0001000010000001: out_v[75] = 10'b1010101000;
    16'b0001100010000000: out_v[75] = 10'b1111010011;
    16'b0000010010000001: out_v[75] = 10'b1000101110;
    16'b0100010010000000: out_v[75] = 10'b1000111010;
    16'b0000000010000001: out_v[75] = 10'b0100101101;
    16'b0010100010010001: out_v[75] = 10'b1000101000;
    16'b0000000010010001: out_v[75] = 10'b0111100011;
    16'b0000010010010001: out_v[75] = 10'b1001011101;
    16'b0010100010000001: out_v[75] = 10'b0110111010;
    16'b0010000000000001: out_v[75] = 10'b0111011110;
    16'b0010000010010000: out_v[75] = 10'b1101001010;
    16'b0010000010000000: out_v[75] = 10'b0111101010;
    16'b0011010010011001: out_v[75] = 10'b1010001011;
    16'b0001000000000001: out_v[75] = 10'b0010111010;
    16'b0001010010011000: out_v[75] = 10'b1101100011;
    16'b0001000010011000: out_v[75] = 10'b0111001011;
    16'b0010010010010000: out_v[75] = 10'b0111110001;
    16'b0010010010000000: out_v[75] = 10'b1111001100;
    16'b0011000010000000: out_v[75] = 10'b1101001001;
    default: out_v[75] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000100100000110: out_v[76] = 10'b0111001011;
    16'b0000101100010010: out_v[76] = 10'b0101100110;
    16'b0000001100010101: out_v[76] = 10'b0100010001;
    16'b0000000100000101: out_v[76] = 10'b0110100011;
    16'b0000000100000010: out_v[76] = 10'b1100001101;
    16'b0000001100000101: out_v[76] = 10'b0110011001;
    16'b0000001100010001: out_v[76] = 10'b1110111111;
    16'b0000000100010101: out_v[76] = 10'b1110011111;
    16'b0000100100000010: out_v[76] = 10'b0011000101;
    16'b0000001100010000: out_v[76] = 10'b1101010001;
    16'b0000101100010000: out_v[76] = 10'b0010100001;
    16'b0000101100010101: out_v[76] = 10'b0110010011;
    16'b0000000100010111: out_v[76] = 10'b0010110100;
    16'b0000001100010111: out_v[76] = 10'b0010101001;
    16'b0000101100010011: out_v[76] = 10'b1111001111;
    16'b0000001100010010: out_v[76] = 10'b1101010001;
    16'b0000100100000111: out_v[76] = 10'b0000100011;
    16'b0000101000010010: out_v[76] = 10'b0000000001;
    16'b0010101100010010: out_v[76] = 10'b0110011110;
    16'b0000100000000010: out_v[76] = 10'b0010001011;
    16'b0000000100000111: out_v[76] = 10'b0010010101;
    16'b0000001000010101: out_v[76] = 10'b1000011101;
    16'b0000100100010010: out_v[76] = 10'b1011101001;
    16'b0000101100000010: out_v[76] = 10'b0110110111;
    16'b0000101100010001: out_v[76] = 10'b0101011111;
    16'b0000001100000111: out_v[76] = 10'b0110100110;
    16'b0000001100010011: out_v[76] = 10'b1001101100;
    16'b0000100100010000: out_v[76] = 10'b1110110111;
    16'b0000000000000101: out_v[76] = 10'b0110010101;
    16'b0000100100000000: out_v[76] = 10'b1111011000;
    16'b0000001000110101: out_v[76] = 10'b1011000110;
    16'b0000101100010111: out_v[76] = 10'b0111011011;
    16'b0000100100000101: out_v[76] = 10'b1001000100;
    16'b0000100100010101: out_v[76] = 10'b0000111011;
    16'b0000100100010111: out_v[76] = 10'b1011011011;
    16'b0000000100000000: out_v[76] = 10'b1001011101;
    16'b0000000001001000: out_v[76] = 10'b0111000111;
    16'b0000000101001000: out_v[76] = 10'b1100000011;
    16'b0010000001001000: out_v[76] = 10'b1111000011;
    16'b0000000000001000: out_v[76] = 10'b1010000110;
    16'b0000100101001000: out_v[76] = 10'b1000001010;
    16'b0000100001001000: out_v[76] = 10'b1000010100;
    16'b0000000101001100: out_v[76] = 10'b1000001111;
    16'b0100000001001000: out_v[76] = 10'b0110001011;
    16'b0100000001001010: out_v[76] = 10'b1010111101;
    16'b0000000101001010: out_v[76] = 10'b1101001100;
    16'b0000000101001101: out_v[76] = 10'b1001111111;
    16'b0000001001001010: out_v[76] = 10'b0010101011;
    16'b0000001001011010: out_v[76] = 10'b1011011110;
    16'b0000000100001000: out_v[76] = 10'b0011101100;
    16'b0000000101001111: out_v[76] = 10'b0011101110;
    16'b0000001101001010: out_v[76] = 10'b1110010011;
    16'b0000001001001000: out_v[76] = 10'b0001100101;
    16'b0000000001001010: out_v[76] = 10'b0111011101;
    16'b0000101001001010: out_v[76] = 10'b0101010100;
    16'b0000001001001110: out_v[76] = 10'b1101000011;
    16'b0000010001001101: out_v[76] = 10'b0111110011;
    16'b0000001001011111: out_v[76] = 10'b1000110111;
    16'b0100001001001010: out_v[76] = 10'b1101001011;
    16'b0000000001001110: out_v[76] = 10'b0010100011;
    16'b0000000101000010: out_v[76] = 10'b1101001010;
    16'b0000000001001111: out_v[76] = 10'b1111000010;
    16'b0100000101001000: out_v[76] = 10'b0110110010;
    16'b0000000001001101: out_v[76] = 10'b0011011000;
    16'b0000001001001111: out_v[76] = 10'b0110010111;
    16'b0000000101001110: out_v[76] = 10'b0110001111;
    16'b0000000100001101: out_v[76] = 10'b1001111110;
    16'b0000100001001010: out_v[76] = 10'b0001110001;
    16'b0000000001001100: out_v[76] = 10'b0111100001;
    16'b0000100100001010: out_v[76] = 10'b0001011101;
    16'b0000100101001110: out_v[76] = 10'b0110111010;
    16'b0000100100001110: out_v[76] = 10'b1000000011;
    16'b0000100000101010: out_v[76] = 10'b0101110111;
    16'b0000000100001010: out_v[76] = 10'b1100000110;
    16'b0000100100001111: out_v[76] = 10'b1100100001;
    16'b0000100000001010: out_v[76] = 10'b1111110010;
    16'b0000000100000110: out_v[76] = 10'b0110100100;
    16'b0000100101001100: out_v[76] = 10'b0110111010;
    16'b0000000000000010: out_v[76] = 10'b0010011011;
    16'b0000100000100010: out_v[76] = 10'b1110101111;
    16'b0000100100001000: out_v[76] = 10'b1100111010;
    16'b0000100101001010: out_v[76] = 10'b0001111000;
    16'b0000000100001111: out_v[76] = 10'b0011011010;
    16'b0000001100000010: out_v[76] = 10'b1101010011;
    16'b0000100101001111: out_v[76] = 10'b1101110010;
    16'b0000100101001101: out_v[76] = 10'b0110001011;
    16'b0000000100001110: out_v[76] = 10'b0100111001;
    16'b0000100001101111: out_v[76] = 10'b0011011111;
    16'b0000000001101111: out_v[76] = 10'b1101001000;
    16'b0000100000101111: out_v[76] = 10'b0000110110;
    16'b0000100001011010: out_v[76] = 10'b1010111010;
    16'b0000001001001011: out_v[76] = 10'b1110010010;
    16'b0000000101001011: out_v[76] = 10'b1011101001;
    16'b0000000001001011: out_v[76] = 10'b0000011101;
    16'b0000100001001111: out_v[76] = 10'b1100110110;
    16'b0000000001101011: out_v[76] = 10'b1111110011;
    16'b0000100101011111: out_v[76] = 10'b0101000010;
    16'b0000100101101111: out_v[76] = 10'b0011011011;
    16'b0000001101001111: out_v[76] = 10'b0110111000;
    16'b0000101101001010: out_v[76] = 10'b0101010110;
    16'b0000100101001011: out_v[76] = 10'b1010010110;
    16'b0000000101011111: out_v[76] = 10'b1110100010;
    16'b0000000101101111: out_v[76] = 10'b0011101111;
    16'b0000101101001111: out_v[76] = 10'b0110110110;
    16'b0000000001101010: out_v[76] = 10'b1011010111;
    16'b0000001101011111: out_v[76] = 10'b1111000011;
    16'b0000100001011000: out_v[76] = 10'b1000101100;
    16'b0000100000000000: out_v[76] = 10'b0000101101;
    16'b0000100101001001: out_v[76] = 10'b1101110000;
    16'b0000101001011000: out_v[76] = 10'b1111000101;
    16'b0000100000001111: out_v[76] = 10'b0101010010;
    16'b0010100100000010: out_v[76] = 10'b1000110111;
    16'b0000100000000111: out_v[76] = 10'b0000011101;
    16'b0000100000100111: out_v[76] = 10'b0101110110;
    16'b0000100101011000: out_v[76] = 10'b0110100111;
    16'b0000100100001011: out_v[76] = 10'b1101100011;
    16'b0010100100001111: out_v[76] = 10'b0010111111;
    16'b0000100000010000: out_v[76] = 10'b1000100111;
    16'b0000100100000011: out_v[76] = 10'b1001001111;
    16'b0010100100001010: out_v[76] = 10'b1100110010;
    16'b0010100100000111: out_v[76] = 10'b1010001110;
    16'b0010100101001000: out_v[76] = 10'b1001001011;
    16'b0100100101001010: out_v[76] = 10'b0000110001;
    16'b1000000101001111: out_v[76] = 10'b1110111111;
    16'b0100100101000010: out_v[76] = 10'b0100010111;
    16'b0100000101001111: out_v[76] = 10'b1111001111;
    16'b1000100101001111: out_v[76] = 10'b1011011110;
    16'b0100100001001010: out_v[76] = 10'b1110101101;
    16'b0010100101001010: out_v[76] = 10'b1101001101;
    16'b0100001101001111: out_v[76] = 10'b1111010001;
    16'b0100100100001010: out_v[76] = 10'b0011111010;
    16'b0100100100000010: out_v[76] = 10'b1110011010;
    16'b0100100100001000: out_v[76] = 10'b1011111111;
    16'b0100100100000000: out_v[76] = 10'b0010100110;
    16'b0100101101001010: out_v[76] = 10'b0101111110;
    16'b0100100101001111: out_v[76] = 10'b1100011011;
    16'b0100100101001000: out_v[76] = 10'b1101101001;
    16'b1000000101001101: out_v[76] = 10'b0100101111;
    16'b0000100101000010: out_v[76] = 10'b0000010111;
    16'b0100000101001010: out_v[76] = 10'b0110111001;
    16'b0000000001011111: out_v[76] = 10'b1010011011;
    16'b0000000100000011: out_v[76] = 10'b0000011011;
    16'b0000000000000011: out_v[76] = 10'b0101110110;
    16'b0000000000100111: out_v[76] = 10'b0111010110;
    16'b0000000001001001: out_v[76] = 10'b0010110101;
    16'b0000000000000111: out_v[76] = 10'b0000111111;
    16'b0000000101001001: out_v[76] = 10'b0010010000;
    16'b0000000101000111: out_v[76] = 10'b0000111101;
    16'b0000000000100011: out_v[76] = 10'b0110000011;
    16'b0000000100100111: out_v[76] = 10'b0111110010;
    16'b0000000100000001: out_v[76] = 10'b0010111011;
    16'b0000000001010111: out_v[76] = 10'b0011101011;
    16'b0000000001000111: out_v[76] = 10'b1000001111;
    16'b0000000000010111: out_v[76] = 10'b0111110000;
    16'b0000000001011011: out_v[76] = 10'b0100011110;
    16'b0000000100010011: out_v[76] = 10'b1001011110;
    16'b0000000000010011: out_v[76] = 10'b1011011011;
    16'b0000100101011101: out_v[76] = 10'b0010101101;
    16'b0000000101011101: out_v[76] = 10'b0100001001;
    16'b0000000001011000: out_v[76] = 10'b0101001110;
    16'b0000100001001101: out_v[76] = 10'b1101000111;
    16'b0000100001101101: out_v[76] = 10'b0101100011;
    16'b0000100001011111: out_v[76] = 10'b1000111010;
    16'b0000100101101101: out_v[76] = 10'b0100110001;
    16'b0000100101011001: out_v[76] = 10'b0111011010;
    16'b0000100100001101: out_v[76] = 10'b0110011111;
    16'b0000000101011000: out_v[76] = 10'b0111010111;
    16'b0000000100001011: out_v[76] = 10'b0000011110;
    16'b0000000000101111: out_v[76] = 10'b1101001011;
    16'b0000000001011010: out_v[76] = 10'b1010101010;
    16'b0000000001100111: out_v[76] = 10'b1010101101;
    16'b0000000100101111: out_v[76] = 10'b1111000000;
    16'b0000001001101111: out_v[76] = 10'b0011110111;
    16'b0000000000001010: out_v[76] = 10'b0101011110;
    default: out_v[76] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000101000000100: out_v[77] = 10'b1010110011;
    16'b0001101000000011: out_v[77] = 10'b1011001011;
    16'b0100101000000011: out_v[77] = 10'b1001011000;
    16'b0001101000000110: out_v[77] = 10'b1011111011;
    16'b0000101000000011: out_v[77] = 10'b0111010010;
    16'b0100100000000001: out_v[77] = 10'b1011001011;
    16'b0010101000000100: out_v[77] = 10'b0101110000;
    16'b0001001000000100: out_v[77] = 10'b1001100001;
    16'b0011101000000011: out_v[77] = 10'b0100011001;
    16'b0011101000000100: out_v[77] = 10'b1000000110;
    16'b0000101000000110: out_v[77] = 10'b0110010101;
    16'b0000101000000101: out_v[77] = 10'b1001100011;
    16'b0011101000000000: out_v[77] = 10'b0011001001;
    16'b0000101000000000: out_v[77] = 10'b0011001101;
    16'b0000100000000011: out_v[77] = 10'b0101111010;
    16'b0001101000000100: out_v[77] = 10'b1011100000;
    16'b0111101000000011: out_v[77] = 10'b0001111011;
    16'b0000000000000011: out_v[77] = 10'b1001001011;
    16'b0100100000000011: out_v[77] = 10'b0011000110;
    16'b0100101000000001: out_v[77] = 10'b1011001011;
    16'b0000100000000000: out_v[77] = 10'b1000001011;
    16'b0001101000000111: out_v[77] = 10'b1011111010;
    16'b0100101000000000: out_v[77] = 10'b0011010011;
    16'b0100000000000011: out_v[77] = 10'b1011010101;
    16'b0001101000000010: out_v[77] = 10'b1001000011;
    16'b0011101000000111: out_v[77] = 10'b1110010011;
    16'b0000101000000010: out_v[77] = 10'b1111010001;
    16'b0011001000000100: out_v[77] = 10'b0111010001;
    16'b0000101000000111: out_v[77] = 10'b1101100011;
    16'b1100000000000011: out_v[77] = 10'b0110011001;
    16'b0101101000000011: out_v[77] = 10'b1111010000;
    16'b0011101000000110: out_v[77] = 10'b0011010101;
    16'b0101000000000011: out_v[77] = 10'b1001000111;
    16'b0001101000000000: out_v[77] = 10'b1101101110;
    16'b0000000000000100: out_v[77] = 10'b0011110011;
    16'b0000100000000010: out_v[77] = 10'b1111010011;
    16'b0000101000000001: out_v[77] = 10'b1110111011;
    16'b0000001000000100: out_v[77] = 10'b1100110011;
    16'b1100000000000001: out_v[77] = 10'b1011001011;
    16'b0100100000000000: out_v[77] = 10'b0011011010;
    16'b0100101000000100: out_v[77] = 10'b0001110101;
    16'b0011000000000000: out_v[77] = 10'b0010001010;
    16'b0000000000000000: out_v[77] = 10'b0010001110;
    16'b0010000000000000: out_v[77] = 10'b0100110001;
    16'b0001000000000000: out_v[77] = 10'b0001111000;
    16'b0011000000000100: out_v[77] = 10'b0010011011;
    16'b1111000000000000: out_v[77] = 10'b1000100111;
    16'b0111000000000000: out_v[77] = 10'b0001010101;
    16'b0110000000000000: out_v[77] = 10'b1000011101;
    16'b0100000000000000: out_v[77] = 10'b1010000011;
    16'b1010000000000000: out_v[77] = 10'b0010001011;
    16'b1100000000000000: out_v[77] = 10'b1001011100;
    16'b0110000000000100: out_v[77] = 10'b0100111101;
    16'b0100000000000010: out_v[77] = 10'b1100110100;
    16'b1111000000000100: out_v[77] = 10'b0001001000;
    16'b0000000000000010: out_v[77] = 10'b1001001110;
    16'b0100000000000110: out_v[77] = 10'b0101100111;
    16'b1000000000000000: out_v[77] = 10'b0110011100;
    16'b0011000000000001: out_v[77] = 10'b0010100100;
    16'b1011000000000000: out_v[77] = 10'b1111010000;
    16'b1110000000000000: out_v[77] = 10'b1010101100;
    16'b0000000000000001: out_v[77] = 10'b0011110110;
    16'b0000000000000110: out_v[77] = 10'b0110010110;
    16'b0110000000000010: out_v[77] = 10'b1011011011;
    16'b0111000000000100: out_v[77] = 10'b0010011110;
    16'b0010000000000010: out_v[77] = 10'b1011001010;
    16'b0100000000000100: out_v[77] = 10'b0111110011;
    16'b0010000000000100: out_v[77] = 10'b0110011000;
    16'b1011000000000001: out_v[77] = 10'b1101000010;
    16'b1011000000000100: out_v[77] = 10'b0010101101;
    16'b1010001000000100: out_v[77] = 10'b0011111110;
    16'b1011101000000100: out_v[77] = 10'b0101010111;
    16'b1011001000000100: out_v[77] = 10'b0110010111;
    16'b0010001000000100: out_v[77] = 10'b1111110000;
    16'b1110000000000100: out_v[77] = 10'b1011101001;
    16'b1111001000000100: out_v[77] = 10'b1000001000;
    16'b1111101000000100: out_v[77] = 10'b0110011010;
    16'b0111001000000100: out_v[77] = 10'b0101001011;
    16'b0010000000000110: out_v[77] = 10'b1011111001;
    16'b1110001000000100: out_v[77] = 10'b0111001011;
    16'b1010000000000100: out_v[77] = 10'b1001000101;
    16'b1110101000000100: out_v[77] = 10'b0111110010;
    16'b1100101000000100: out_v[77] = 10'b1110000100;
    16'b0111101000000100: out_v[77] = 10'b1100000111;
    16'b0110101000000100: out_v[77] = 10'b0111110110;
    16'b0011000000000010: out_v[77] = 10'b1010101110;
    16'b1111101000000101: out_v[77] = 10'b0100011011;
    16'b0110001000000100: out_v[77] = 10'b0101101011;
    16'b0011100000000000: out_v[77] = 10'b0000110111;
    16'b0010101000000101: out_v[77] = 10'b1001111010;
    16'b0000101001000100: out_v[77] = 10'b1010001111;
    16'b0010100000000000: out_v[77] = 10'b1100100001;
    16'b0010101000000000: out_v[77] = 10'b0111111001;
    16'b0010101000000110: out_v[77] = 10'b1110101010;
    16'b0010101000000011: out_v[77] = 10'b1110001011;
    16'b0010101000000010: out_v[77] = 10'b1001100001;
    16'b0011101000000101: out_v[77] = 10'b0100011111;
    16'b1100000000000010: out_v[77] = 10'b0011010011;
    16'b0010101000000111: out_v[77] = 10'b1000100010;
    16'b0001000000000100: out_v[77] = 10'b1011100100;
    16'b0100001000000100: out_v[77] = 10'b1111000010;
    16'b0011101001000100: out_v[77] = 10'b0010101010;
    16'b0001101001000100: out_v[77] = 10'b1000010111;
    16'b0001001001000100: out_v[77] = 10'b1011001011;
    16'b1110101000000101: out_v[77] = 10'b1111110010;
    16'b0000101001000000: out_v[77] = 10'b0101110100;
    16'b0101101000000100: out_v[77] = 10'b0100100010;
    16'b0000101010000100: out_v[77] = 10'b0100000111;
    16'b0000001010000100: out_v[77] = 10'b1010101100;
    16'b0010101000000001: out_v[77] = 10'b0110101010;
    16'b0000100000000001: out_v[77] = 10'b0011111110;
    16'b0000000010000100: out_v[77] = 10'b0111011001;
    16'b0110101000000101: out_v[77] = 10'b1111010110;
    16'b0000101010000101: out_v[77] = 10'b1110111011;
    16'b0100101000000101: out_v[77] = 10'b1011001001;
    16'b0000101010000000: out_v[77] = 10'b0001001001;
    16'b1001000000000000: out_v[77] = 10'b1101100111;
    16'b0001100000000000: out_v[77] = 10'b0011110110;
    16'b1011101000000000: out_v[77] = 10'b0011011111;
    16'b0011001000000000: out_v[77] = 10'b1011101011;
    16'b1010101000000100: out_v[77] = 10'b1100111110;
    16'b0010001000000000: out_v[77] = 10'b1011100010;
    16'b1000101000000100: out_v[77] = 10'b0110100011;
    16'b0010100000000100: out_v[77] = 10'b1101100011;
    16'b0011100000000100: out_v[77] = 10'b0101000111;
    16'b0111101000000000: out_v[77] = 10'b0111001111;
    default: out_v[77] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000000010000: out_v[78] = 10'b0100101101;
    16'b0000000000110000: out_v[78] = 10'b1001100101;
    16'b0000001000100100: out_v[78] = 10'b0110011011;
    16'b0000101000100000: out_v[78] = 10'b1110001001;
    16'b0000000000000000: out_v[78] = 10'b0000101010;
    16'b0000101000000100: out_v[78] = 10'b1010100010;
    16'b0000000000100000: out_v[78] = 10'b1010001101;
    16'b0000001000000000: out_v[78] = 10'b0101111000;
    16'b0000001000100000: out_v[78] = 10'b0100000001;
    16'b0000001000110000: out_v[78] = 10'b1000010101;
    16'b0000000010010000: out_v[78] = 10'b1100111110;
    16'b0000101000100100: out_v[78] = 10'b0001010011;
    16'b0000100000100100: out_v[78] = 10'b1011001001;
    16'b0000001000000100: out_v[78] = 10'b1011100110;
    16'b0000001000010000: out_v[78] = 10'b0101100100;
    16'b0000000000100100: out_v[78] = 10'b0011000100;
    16'b0000000010000000: out_v[78] = 10'b1000110010;
    16'b0000000010110000: out_v[78] = 10'b0100100010;
    16'b0000001010010000: out_v[78] = 10'b0101111000;
    16'b0000001010000000: out_v[78] = 10'b0001011110;
    16'b0000000000010100: out_v[78] = 10'b1100001100;
    16'b0000001010110000: out_v[78] = 10'b1000011110;
    16'b0000000010100000: out_v[78] = 10'b0110010110;
    16'b0000000000000100: out_v[78] = 10'b0110010101;
    16'b0000000010000100: out_v[78] = 10'b0010010110;
    16'b0000001000010100: out_v[78] = 10'b1010101111;
    16'b0000001010000100: out_v[78] = 10'b0000111010;
    16'b0001001000010000: out_v[78] = 10'b1011000110;
    16'b0000000010010100: out_v[78] = 10'b0110001010;
    16'b0001001010010000: out_v[78] = 10'b0011100101;
    16'b0000001010010100: out_v[78] = 10'b0010001100;
    16'b0001000000010000: out_v[78] = 10'b1010110110;
    16'b0000001010100000: out_v[78] = 10'b1110111001;
    16'b0000000010110100: out_v[78] = 10'b0100111010;
    16'b0000100010110100: out_v[78] = 10'b1100110010;
    16'b0000101010110100: out_v[78] = 10'b1110110010;
    16'b0000100000110100: out_v[78] = 10'b1101110111;
    16'b0000101010010100: out_v[78] = 10'b0100111010;
    16'b0000100010010100: out_v[78] = 10'b1001110001;
    16'b0010001010010000: out_v[78] = 10'b1111010011;
    16'b0010001010000000: out_v[78] = 10'b0010101111;
    16'b0010001000010000: out_v[78] = 10'b0110011111;
    16'b0000000010100100: out_v[78] = 10'b0110010010;
    16'b0000100010100100: out_v[78] = 10'b0111110101;
    16'b0000100000100000: out_v[78] = 10'b0110000110;
    16'b0000100000000100: out_v[78] = 10'b0011100011;
    16'b0000001010110100: out_v[78] = 10'b0110000100;
    16'b0000000000110100: out_v[78] = 10'b1110100010;
    default: out_v[78] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1000000001101011: out_v[79] = 10'b0110100000;
    16'b1000000001101001: out_v[79] = 10'b0001001011;
    16'b1000000001101000: out_v[79] = 10'b1110010101;
    16'b0000000001101010: out_v[79] = 10'b1000101101;
    16'b1000000000100010: out_v[79] = 10'b0000101111;
    16'b1000001001101001: out_v[79] = 10'b1010100110;
    16'b0000000001001000: out_v[79] = 10'b0000111011;
    16'b1000001001001001: out_v[79] = 10'b1001000110;
    16'b0000000000001000: out_v[79] = 10'b0001101001;
    16'b0000000001100010: out_v[79] = 10'b0010010101;
    16'b1000000001101010: out_v[79] = 10'b0001011111;
    16'b0000000001101000: out_v[79] = 10'b1010000101;
    16'b1000000001100010: out_v[79] = 10'b1010001110;
    16'b0000000001001010: out_v[79] = 10'b1111010110;
    16'b1000000001100011: out_v[79] = 10'b1101001011;
    16'b1000000001001010: out_v[79] = 10'b0110011011;
    16'b1000000001000011: out_v[79] = 10'b1100100001;
    16'b1000000000101001: out_v[79] = 10'b1010101100;
    16'b0000000000101000: out_v[79] = 10'b1101101101;
    16'b1000000001001011: out_v[79] = 10'b0100011001;
    16'b0000000001000010: out_v[79] = 10'b0000100011;
    16'b1000001001101011: out_v[79] = 10'b0000001011;
    16'b0000000000100010: out_v[79] = 10'b0000011101;
    16'b1000000001001000: out_v[79] = 10'b1101101000;
    16'b0000000001100000: out_v[79] = 10'b1110100111;
    16'b1000000001000010: out_v[79] = 10'b1011101001;
    16'b1000000000000011: out_v[79] = 10'b1010100100;
    16'b1000001011101011: out_v[79] = 10'b1101010110;
    16'b1000000000101000: out_v[79] = 10'b1011111110;
    16'b0000000000000010: out_v[79] = 10'b1010100011;
    16'b1000000001001001: out_v[79] = 10'b0111100001;
    16'b1000001011101001: out_v[79] = 10'b1000100100;
    16'b0000000000101010: out_v[79] = 10'b1001011101;
    16'b1000001001101000: out_v[79] = 10'b1101001011;
    16'b1000000000101011: out_v[79] = 10'b1011000011;
    16'b1000000000001011: out_v[79] = 10'b1000011111;
    16'b0000000011100000: out_v[79] = 10'b0010101011;
    16'b0000001010100000: out_v[79] = 10'b0101100111;
    16'b0000001010001000: out_v[79] = 10'b0101111100;
    16'b0000001010001010: out_v[79] = 10'b0001111010;
    16'b0000000010000000: out_v[79] = 10'b1101011011;
    16'b0000000010001010: out_v[79] = 10'b0101000010;
    16'b0000000011000000: out_v[79] = 10'b1110100011;
    16'b0000001000001010: out_v[79] = 10'b0101010010;
    16'b0000001011100000: out_v[79] = 10'b0000110010;
    16'b0000001010000000: out_v[79] = 10'b0001111110;
    16'b0000001011000000: out_v[79] = 10'b0000111001;
    16'b0000000010001000: out_v[79] = 10'b1100001111;
    16'b0000001011101000: out_v[79] = 10'b1010001100;
    16'b0000000010100000: out_v[79] = 10'b1001100011;
    16'b0000001010000010: out_v[79] = 10'b0100100101;
    16'b0000001010101000: out_v[79] = 10'b0011100110;
    16'b0000001000001000: out_v[79] = 10'b1100100110;
    16'b0000001011001000: out_v[79] = 10'b0011100111;
    16'b0000001011001010: out_v[79] = 10'b0100000100;
    16'b1000001001100011: out_v[79] = 10'b0011100110;
    16'b0000001011000010: out_v[79] = 10'b0001000100;
    16'b0000000011100010: out_v[79] = 10'b0001110101;
    16'b0000001011100010: out_v[79] = 10'b0110101011;
    16'b1000001011000011: out_v[79] = 10'b1100011100;
    16'b0000001010000011: out_v[79] = 10'b1111100010;
    16'b1000001011100011: out_v[79] = 10'b0010101011;
    16'b0000000010000010: out_v[79] = 10'b0011101100;
    16'b0000001011100011: out_v[79] = 10'b0000110111;
    16'b1000001010100011: out_v[79] = 10'b0100110010;
    16'b0000000011000010: out_v[79] = 10'b1001110100;
    16'b0000001011000011: out_v[79] = 10'b1001101111;
    16'b0000001010100010: out_v[79] = 10'b1111001000;
    16'b1000001010101001: out_v[79] = 10'b1011110010;
    16'b1000001010000011: out_v[79] = 10'b1111000001;
    16'b0000001011001011: out_v[79] = 10'b1000001110;
    16'b1000001001000011: out_v[79] = 10'b1011000111;
    16'b0000001001000011: out_v[79] = 10'b0011110100;
    16'b0000001011101011: out_v[79] = 10'b0001110111;
    16'b1000001010001001: out_v[79] = 10'b0010100101;
    16'b0000001011101010: out_v[79] = 10'b1001100001;
    16'b0000001011101001: out_v[79] = 10'b0010100111;
    16'b1000001011001011: out_v[79] = 10'b0011011010;
    16'b1000001011100001: out_v[79] = 10'b0101011100;
    16'b1000001011001001: out_v[79] = 10'b0111000110;
    16'b1000001010100001: out_v[79] = 10'b1000110010;
    16'b0000000000000011: out_v[79] = 10'b1001101011;
    16'b0000000001100011: out_v[79] = 10'b1101001010;
    16'b1000000000000001: out_v[79] = 10'b0010110000;
    16'b1000000000100011: out_v[79] = 10'b0100100011;
    16'b0000001000000000: out_v[79] = 10'b1001010000;
    16'b0000001000000010: out_v[79] = 10'b1001100001;
    16'b0000000001000011: out_v[79] = 10'b0111111011;
    16'b1000001001001011: out_v[79] = 10'b0110001110;
    16'b0000001001100010: out_v[79] = 10'b0111010010;
    16'b0000001001100011: out_v[79] = 10'b0101011011;
    16'b1000000000001001: out_v[79] = 10'b1011100110;
    16'b0000001000100010: out_v[79] = 10'b0111001111;
    16'b0000000000100011: out_v[79] = 10'b0111011111;
    16'b1000000000100001: out_v[79] = 10'b0101011110;
    16'b1000000001100001: out_v[79] = 10'b1001011010;
    16'b0000001001000010: out_v[79] = 10'b0010011010;
    16'b0000000000001011: out_v[79] = 10'b0010011011;
    16'b0000001010000001: out_v[79] = 10'b0101110011;
    16'b1000001010000001: out_v[79] = 10'b0100011101;
    16'b0000001000001001: out_v[79] = 10'b1111000010;
    16'b1000001000000001: out_v[79] = 10'b0000010010;
    16'b0000000000000001: out_v[79] = 10'b1011011111;
    16'b1000001000001011: out_v[79] = 10'b1010110101;
    16'b1000001000100001: out_v[79] = 10'b1101011000;
    16'b1000001010101011: out_v[79] = 10'b1101011000;
    16'b0000001000100000: out_v[79] = 10'b0111000110;
    16'b0000001010101001: out_v[79] = 10'b1001001010;
    16'b0000001000100001: out_v[79] = 10'b0111001011;
    16'b0000001000000001: out_v[79] = 10'b0101110001;
    16'b0000001010100001: out_v[79] = 10'b0010110100;
    16'b1000000010000001: out_v[79] = 10'b0011100111;
    16'b0000001000101000: out_v[79] = 10'b0110010000;
    16'b0000001010001001: out_v[79] = 10'b1000011000;
    16'b1000001010001011: out_v[79] = 10'b0111010000;
    16'b1000001000001001: out_v[79] = 10'b1100100011;
    16'b1000001000101001: out_v[79] = 10'b0010100001;
    16'b1000000010100001: out_v[79] = 10'b1001011101;
    16'b0000001000101001: out_v[79] = 10'b1101010111;
    16'b1010001010001001: out_v[79] = 10'b0111000100;
    16'b1010001010000001: out_v[79] = 10'b1110001010;
    16'b0000001010001011: out_v[79] = 10'b0010011110;
    16'b0000001001000000: out_v[79] = 10'b1101101000;
    16'b0000001001101000: out_v[79] = 10'b0110111001;
    16'b0000000000101001: out_v[79] = 10'b0010111111;
    16'b1010000001101001: out_v[79] = 10'b0111011111;
    16'b0010001011101000: out_v[79] = 10'b0010111010;
    16'b0000000001101001: out_v[79] = 10'b0100011011;
    16'b0000001001101001: out_v[79] = 10'b0010101001;
    16'b0000001001001000: out_v[79] = 10'b1111110011;
    16'b0010001001101000: out_v[79] = 10'b0001011110;
    16'b0010001010101000: out_v[79] = 10'b1111000010;
    16'b1000000000000010: out_v[79] = 10'b1011100011;
    16'b0000001001101010: out_v[79] = 10'b1110101001;
    16'b0000000010101000: out_v[79] = 10'b0001111100;
    16'b0000000001001001: out_v[79] = 10'b1010110110;
    16'b0000000110000010: out_v[79] = 10'b1110111000;
    16'b1000001110001011: out_v[79] = 10'b1101000110;
    16'b1000000110000011: out_v[79] = 10'b1111101110;
    16'b1000000010001011: out_v[79] = 10'b1110010011;
    16'b1000001100001011: out_v[79] = 10'b1111000111;
    16'b1000000010000011: out_v[79] = 10'b0110100111;
    16'b1000000010001001: out_v[79] = 10'b1101001111;
    16'b1000001000000011: out_v[79] = 10'b1010100110;
    16'b1000001111001011: out_v[79] = 10'b1111110011;
    16'b1000001110000011: out_v[79] = 10'b0000111011;
    16'b0000000000001001: out_v[79] = 10'b0011100101;
    16'b1000000011001001: out_v[79] = 10'b1111011010;
    16'b1000000100001011: out_v[79] = 10'b1110101101;
    16'b1000001100000011: out_v[79] = 10'b1110111101;
    16'b1000000110001011: out_v[79] = 10'b1110011011;
    16'b0000000000000000: out_v[79] = 10'b0011101000;
    16'b1000001010000000: out_v[79] = 10'b1001011000;
    16'b1000000010000010: out_v[79] = 10'b1111100100;
    16'b1000000100000011: out_v[79] = 10'b1111110110;
    16'b1001001000001001: out_v[79] = 10'b0001111111;
    16'b1000000000001000: out_v[79] = 10'b0011000101;
    16'b0000000011001000: out_v[79] = 10'b0111011000;
    16'b0000000011101000: out_v[79] = 10'b1001010100;
    16'b0000001010101010: out_v[79] = 10'b0011111011;
    16'b0000000010000011: out_v[79] = 10'b0111010011;
    16'b0000001001001010: out_v[79] = 10'b1110110011;
    16'b0000001000101010: out_v[79] = 10'b0110110100;
    16'b1000000010101001: out_v[79] = 10'b0101011001;
    default: out_v[79] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100010000000000: out_v[80] = 10'b0000100001;
    16'b0001110000000000: out_v[80] = 10'b0011110011;
    16'b0101110000000000: out_v[80] = 10'b0100000001;
    16'b0010110000000000: out_v[80] = 10'b1011110010;
    16'b0011110000000000: out_v[80] = 10'b0011110100;
    16'b0101100000000000: out_v[80] = 10'b0101000001;
    16'b0000110000000000: out_v[80] = 10'b1100011001;
    16'b0111110000000000: out_v[80] = 10'b0001010001;
    16'b0100110000000000: out_v[80] = 10'b0101111000;
    16'b0010100000000000: out_v[80] = 10'b0110010001;
    16'b0110110000000000: out_v[80] = 10'b1001011100;
    16'b0101110001000000: out_v[80] = 10'b1010100011;
    16'b0011100000000000: out_v[80] = 10'b1101100110;
    16'b0110010000000000: out_v[80] = 10'b1110100110;
    16'b0101010000000000: out_v[80] = 10'b1100010111;
    16'b0001100000000000: out_v[80] = 10'b1100011101;
    16'b0001010000000000: out_v[80] = 10'b1011000100;
    16'b0000010000000000: out_v[80] = 10'b0101110010;
    16'b0100100000000000: out_v[80] = 10'b0001000101;
    16'b0111100000000000: out_v[80] = 10'b1100000110;
    16'b0110100000000000: out_v[80] = 10'b1010010111;
    16'b0000100000000000: out_v[80] = 10'b0010100111;
    16'b0101000000000000: out_v[80] = 10'b0010111001;
    16'b0010000000000000: out_v[80] = 10'b0111011000;
    16'b0100000000000000: out_v[80] = 10'b1010001101;
    16'b0110000000000000: out_v[80] = 10'b1010100010;
    16'b0000000000000000: out_v[80] = 10'b0010110010;
    16'b0010010000000000: out_v[80] = 10'b0111110101;
    16'b0110010000000010: out_v[80] = 10'b0010011011;
    16'b0110110000000010: out_v[80] = 10'b1000010110;
    16'b0100000000000010: out_v[80] = 10'b1000001010;
    16'b0100010000000010: out_v[80] = 10'b0101101110;
    16'b0100100000000010: out_v[80] = 10'b1001010111;
    16'b0111000000000000: out_v[80] = 10'b1010010001;
    16'b0011000000000000: out_v[80] = 10'b0010010011;
    16'b0001000000000000: out_v[80] = 10'b0111110000;
    16'b0000010001000000: out_v[80] = 10'b0111010010;
    16'b0111010000000000: out_v[80] = 10'b0001111010;
    16'b0011010000000000: out_v[80] = 10'b1101000101;
    16'b0010000001000000: out_v[80] = 10'b0010110011;
    16'b0010010001000000: out_v[80] = 10'b0110001101;
    16'b0000010001001000: out_v[80] = 10'b1111100111;
    16'b0001010001000000: out_v[80] = 10'b1011001010;
    16'b0011000001000000: out_v[80] = 10'b0010111011;
    16'b0000000001000000: out_v[80] = 10'b1111101001;
    default: out_v[80] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001000000000000: out_v[81] = 10'b0111110011;
    16'b0010000010001000: out_v[81] = 10'b1011100110;
    16'b0110000010001000: out_v[81] = 10'b0010010111;
    16'b0000000000001000: out_v[81] = 10'b0110010111;
    16'b0111010000000000: out_v[81] = 10'b1010100011;
    16'b0101010010001000: out_v[81] = 10'b1000101001;
    16'b0000000010000000: out_v[81] = 10'b0000110011;
    16'b0000000010100010: out_v[81] = 10'b1110011111;
    16'b0011010000000000: out_v[81] = 10'b1000010111;
    16'b0000000010001000: out_v[81] = 10'b1000011101;
    16'b0100000010001000: out_v[81] = 10'b1110000111;
    16'b0000000010001010: out_v[81] = 10'b0100001111;
    16'b0000000000001010: out_v[81] = 10'b0000011001;
    16'b0010000000001010: out_v[81] = 10'b0000110101;
    16'b0110000000001000: out_v[81] = 10'b0101000111;
    16'b0111000000001010: out_v[81] = 10'b1011101010;
    16'b0100000000001010: out_v[81] = 10'b0110011100;
    16'b0011000000001010: out_v[81] = 10'b0010011011;
    16'b0011000000001000: out_v[81] = 10'b1111110000;
    16'b0100000010001010: out_v[81] = 10'b0000000111;
    16'b0000000000101010: out_v[81] = 10'b1010010110;
    16'b0101010000000000: out_v[81] = 10'b0111100001;
    16'b0001000000001010: out_v[81] = 10'b1000101000;
    16'b0111000000001000: out_v[81] = 10'b0001110010;
    16'b0000000001101010: out_v[81] = 10'b1000011101;
    16'b0100000010101010: out_v[81] = 10'b0110110111;
    16'b0100010010001000: out_v[81] = 10'b1110000101;
    16'b0100000010000000: out_v[81] = 10'b0011110101;
    16'b0100000000001000: out_v[81] = 10'b0110100111;
    16'b0001010000000000: out_v[81] = 10'b0111000101;
    16'b0011000010001000: out_v[81] = 10'b1000011011;
    16'b0111010010001000: out_v[81] = 10'b0010011001;
    16'b0000000010000010: out_v[81] = 10'b1010000101;
    16'b0111010000001000: out_v[81] = 10'b1010101010;
    16'b0111010000000010: out_v[81] = 10'b0011010000;
    16'b0011000000000010: out_v[81] = 10'b1100011010;
    16'b0101010010000000: out_v[81] = 10'b1010011111;
    16'b0011000000000000: out_v[81] = 10'b0110010101;
    16'b0111010000001010: out_v[81] = 10'b0010011011;
    16'b0000000010101010: out_v[81] = 10'b1011100101;
    16'b0001000010001000: out_v[81] = 10'b0101110110;
    16'b0011010000000010: out_v[81] = 10'b1001000011;
    16'b0001000000000010: out_v[81] = 10'b0111001001;
    16'b0000000000000000: out_v[81] = 10'b0101001110;
    16'b0110010010001000: out_v[81] = 10'b0000011111;
    16'b0111000010001000: out_v[81] = 10'b1101011011;
    16'b0011000000101010: out_v[81] = 10'b0110101011;
    16'b0010000010001010: out_v[81] = 10'b0101110011;
    16'b0000000000100010: out_v[81] = 10'b1010010101;
    16'b0010000000001000: out_v[81] = 10'b1101000100;
    16'b0111000000000000: out_v[81] = 10'b0100101100;
    16'b0100000000000000: out_v[81] = 10'b1010000110;
    16'b0100000000000010: out_v[81] = 10'b1001000011;
    16'b0010000000000000: out_v[81] = 10'b0111101000;
    16'b0111000010000000: out_v[81] = 10'b0101001110;
    16'b0110000000000000: out_v[81] = 10'b0110100011;
    16'b0011000010000000: out_v[81] = 10'b1001100111;
    16'b0100010000000010: out_v[81] = 10'b0101011111;
    16'b0010000010000000: out_v[81] = 10'b1110101010;
    16'b0000000000000010: out_v[81] = 10'b1010001111;
    16'b0110010000000000: out_v[81] = 10'b0110110011;
    16'b0110000001000010: out_v[81] = 10'b0111000001;
    16'b0110010000000010: out_v[81] = 10'b1110001111;
    16'b0110000000100010: out_v[81] = 10'b0111001101;
    16'b0100000000100000: out_v[81] = 10'b1100000100;
    16'b0011010000100000: out_v[81] = 10'b0101110111;
    16'b0111010000100010: out_v[81] = 10'b1000100110;
    16'b0010000001000010: out_v[81] = 10'b1011000100;
    16'b0010000000000010: out_v[81] = 10'b0111101100;
    16'b0111000000000010: out_v[81] = 10'b0101011001;
    16'b0111010011000010: out_v[81] = 10'b1001000111;
    16'b0101010011001010: out_v[81] = 10'b1110110111;
    16'b0100010010001010: out_v[81] = 10'b1010010101;
    16'b0111010000100000: out_v[81] = 10'b0000010100;
    16'b0110000000000010: out_v[81] = 10'b1000111101;
    16'b0101010000000010: out_v[81] = 10'b0001111100;
    16'b0111000000100010: out_v[81] = 10'b1011111101;
    16'b0111010001000010: out_v[81] = 10'b0000000100;
    16'b0110000000100000: out_v[81] = 10'b1011000011;
    16'b0101010000001010: out_v[81] = 10'b0001001111;
    16'b0111010001100010: out_v[81] = 10'b1101110111;
    16'b0101010010000010: out_v[81] = 10'b1000011100;
    16'b0101010001000010: out_v[81] = 10'b1001110100;
    16'b0001010010000000: out_v[81] = 10'b0101011010;
    16'b0111000001000010: out_v[81] = 10'b1011110110;
    16'b0111010010000010: out_v[81] = 10'b1111000001;
    16'b0011010001000010: out_v[81] = 10'b1101011011;
    16'b0011000001000010: out_v[81] = 10'b1001001001;
    16'b0101010000100010: out_v[81] = 10'b1110111001;
    16'b0111010010000000: out_v[81] = 10'b0010011010;
    16'b0100000000100010: out_v[81] = 10'b0110010110;
    16'b0010000000100010: out_v[81] = 10'b0101010100;
    16'b0101010010001010: out_v[81] = 10'b1011110011;
    16'b0101010011000010: out_v[81] = 10'b1111001110;
    16'b0011010000100010: out_v[81] = 10'b1001111110;
    16'b0111000010000010: out_v[81] = 10'b1001001010;
    16'b0010010000000010: out_v[81] = 10'b1111001000;
    16'b0000010000000010: out_v[81] = 10'b1010111100;
    16'b0001010010000010: out_v[81] = 10'b0100011010;
    16'b0001010000000010: out_v[81] = 10'b1100111010;
    16'b0000010001000010: out_v[81] = 10'b1011101000;
    16'b0010010000000000: out_v[81] = 10'b0101011011;
    16'b0011010010000000: out_v[81] = 10'b0010011001;
    16'b0011010010000010: out_v[81] = 10'b0110000000;
    16'b0010010010000010: out_v[81] = 10'b1110001100;
    16'b0010010010000000: out_v[81] = 10'b1101111010;
    16'b0010010001000010: out_v[81] = 10'b0101010010;
    16'b0000010000000000: out_v[81] = 10'b0001111000;
    16'b0011000010000010: out_v[81] = 10'b1001111110;
    16'b0110010000001000: out_v[81] = 10'b1100010110;
    16'b0011010001000000: out_v[81] = 10'b0001010011;
    16'b0011010000001000: out_v[81] = 10'b0010111010;
    16'b0011110000000000: out_v[81] = 10'b0001110111;
    16'b0001010010001000: out_v[81] = 10'b0100011001;
    16'b0101010000001000: out_v[81] = 10'b1001110010;
    16'b0100010000000000: out_v[81] = 10'b0111111000;
    16'b0000010010000010: out_v[81] = 10'b1011110110;
    16'b0100010010000000: out_v[81] = 10'b0010100000;
    16'b0000010010000000: out_v[81] = 10'b0001110100;
    16'b0100010010000010: out_v[81] = 10'b0001100011;
    16'b0110000010000000: out_v[81] = 10'b0011100000;
    16'b0001000010000000: out_v[81] = 10'b0110011000;
    16'b0110010010000000: out_v[81] = 10'b0001101000;
    16'b0001000010000010: out_v[81] = 10'b1011101010;
    16'b0101000000001010: out_v[81] = 10'b0110100010;
    16'b0101010000101000: out_v[81] = 10'b0111101011;
    16'b0100010000101010: out_v[81] = 10'b0011011010;
    16'b0100010000001010: out_v[81] = 10'b0111000000;
    16'b0101000000000010: out_v[81] = 10'b1101001010;
    16'b0101000000001000: out_v[81] = 10'b1111001000;
    16'b0101000000000000: out_v[81] = 10'b0100011001;
    16'b0100010000001000: out_v[81] = 10'b0111010000;
    16'b0101000000101010: out_v[81] = 10'b0011101000;
    16'b0101010000101010: out_v[81] = 10'b1110101000;
    16'b0100010000100010: out_v[81] = 10'b0011101010;
    16'b0111000000101010: out_v[81] = 10'b1110111001;
    16'b0001000000001000: out_v[81] = 10'b0011110110;
    16'b0011110000000001: out_v[81] = 10'b0111011010;
    16'b0111110000000000: out_v[81] = 10'b0011100111;
    16'b0101000010000000: out_v[81] = 10'b1110001000;
    16'b0001010010001010: out_v[81] = 10'b0001111110;
    16'b0101000010000010: out_v[81] = 10'b0110001111;
    16'b0011110000001000: out_v[81] = 10'b0111111010;
    16'b0010110000000000: out_v[81] = 10'b1110001100;
    16'b0001110000000000: out_v[81] = 10'b1001100111;
    16'b0000110000000000: out_v[81] = 10'b1110010001;
    default: out_v[81] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010100000100000: out_v[82] = 10'b1000110111;
    16'b0000000000000000: out_v[82] = 10'b0011110001;
    16'b0010100000000000: out_v[82] = 10'b0000011101;
    16'b0010000000000000: out_v[82] = 10'b1000100101;
    16'b0000100000100000: out_v[82] = 10'b1110010001;
    16'b0000100000000000: out_v[82] = 10'b0111001001;
    16'b0010000010000000: out_v[82] = 10'b1111000101;
    16'b1000100000000000: out_v[82] = 10'b1101101011;
    16'b1000100000100000: out_v[82] = 10'b1000000111;
    16'b0010100010000000: out_v[82] = 10'b0000110111;
    16'b1000000000000000: out_v[82] = 10'b1110101111;
    16'b0010000000100000: out_v[82] = 10'b1101100011;
    16'b1010000000000000: out_v[82] = 10'b1000001101;
    16'b1000000000100000: out_v[82] = 10'b1011100000;
    16'b0000000000100000: out_v[82] = 10'b1111000110;
    16'b1010100000000000: out_v[82] = 10'b1111001010;
    16'b0010100010100000: out_v[82] = 10'b0001010110;
    16'b1010100000100000: out_v[82] = 10'b0001101110;
    16'b1000000000001000: out_v[82] = 10'b1110000010;
    16'b1010000000001000: out_v[82] = 10'b0100010111;
    16'b1000100000001000: out_v[82] = 10'b1100011010;
    16'b1010000010001010: out_v[82] = 10'b1111010000;
    16'b0010100000101000: out_v[82] = 10'b1100011100;
    16'b1010000010001000: out_v[82] = 10'b1000101011;
    16'b0010000000001000: out_v[82] = 10'b0101011100;
    16'b1010100000001000: out_v[82] = 10'b0111111000;
    16'b1010000010001001: out_v[82] = 10'b1101001101;
    16'b0010000000101000: out_v[82] = 10'b1011110110;
    16'b0010000010100000: out_v[82] = 10'b1001000011;
    16'b1000100000101000: out_v[82] = 10'b1001001110;
    16'b0010100010100011: out_v[82] = 10'b1110010111;
    16'b1010100000101000: out_v[82] = 10'b1110000000;
    16'b0000100000001000: out_v[82] = 10'b1101001100;
    16'b0010100010100010: out_v[82] = 10'b1110000100;
    16'b0000100000101000: out_v[82] = 10'b1010001100;
    16'b1010000010001011: out_v[82] = 10'b1101010101;
    16'b1010000000101000: out_v[82] = 10'b0010111111;
    16'b1010100010101000: out_v[82] = 10'b1111001010;
    16'b1010100010001011: out_v[82] = 10'b0100011111;
    16'b1010100010001000: out_v[82] = 10'b1111000110;
    16'b0010100010100001: out_v[82] = 10'b0001110111;
    16'b0010110010100011: out_v[82] = 10'b1100101111;
    16'b1010000010000010: out_v[82] = 10'b1011001101;
    16'b0010100000001000: out_v[82] = 10'b0101101110;
    16'b0010100010101000: out_v[82] = 10'b1011001101;
    16'b1010010010001011: out_v[82] = 10'b1111010111;
    16'b1010000010101000: out_v[82] = 10'b0011101001;
    16'b1010000010000000: out_v[82] = 10'b1111001101;
    16'b0010100010001000: out_v[82] = 10'b1111110010;
    16'b1000000000101000: out_v[82] = 10'b0000111100;
    16'b1010000000100000: out_v[82] = 10'b0111111010;
    16'b1010000010101011: out_v[82] = 10'b1111010110;
    16'b1010000010101001: out_v[82] = 10'b0011001011;
    16'b1010000010100000: out_v[82] = 10'b1110000011;
    16'b1010000010101010: out_v[82] = 10'b0010110011;
    16'b0010000010101000: out_v[82] = 10'b0010100110;
    16'b1010000010100001: out_v[82] = 10'b1100010100;
    16'b1010010010101011: out_v[82] = 10'b1010001000;
    16'b1010100010000000: out_v[82] = 10'b0111110010;
    16'b1010000010100010: out_v[82] = 10'b0011011011;
    16'b1010100010101010: out_v[82] = 10'b1110110110;
    16'b1010100010101001: out_v[82] = 10'b0101001010;
    16'b1010100010101011: out_v[82] = 10'b0101101110;
    16'b1010111010101011: out_v[82] = 10'b0100110111;
    16'b1010011010101011: out_v[82] = 10'b0011101110;
    16'b1010000010100011: out_v[82] = 10'b1110100010;
    16'b1010100010100000: out_v[82] = 10'b0100100110;
    16'b0000000000101000: out_v[82] = 10'b1111100100;
    16'b0000100010100010: out_v[82] = 10'b1100110011;
    16'b0000100010101000: out_v[82] = 10'b0010111011;
    16'b1000000010101000: out_v[82] = 10'b0000011010;
    16'b0000000000001000: out_v[82] = 10'b0010111000;
    16'b1000100010101000: out_v[82] = 10'b0111010110;
    16'b0000100010100000: out_v[82] = 10'b0110000011;
    16'b0000100010100011: out_v[82] = 10'b0100111010;
    16'b0000000010100000: out_v[82] = 10'b0110110010;
    16'b0000100000100001: out_v[82] = 10'b0101011110;
    16'b1000000000001001: out_v[82] = 10'b0111110101;
    16'b1000000010001000: out_v[82] = 10'b1101010101;
    16'b0000101000100001: out_v[82] = 10'b1000110000;
    16'b0000100010100001: out_v[82] = 10'b1101000110;
    16'b0000100000101001: out_v[82] = 10'b1111101001;
    16'b1000100000101001: out_v[82] = 10'b0010001111;
    16'b0000000000100001: out_v[82] = 10'b0011110111;
    default: out_v[82] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100100011010000: out_v[83] = 10'b0001010111;
    16'b0010000011010000: out_v[83] = 10'b1001011010;
    16'b0000001011010000: out_v[83] = 10'b0000100010;
    16'b0100000011010000: out_v[83] = 10'b0100100100;
    16'b0000000001000000: out_v[83] = 10'b1011101011;
    16'b0010000011000000: out_v[83] = 10'b0010001011;
    16'b0000001001000000: out_v[83] = 10'b1000110001;
    16'b0000000001010000: out_v[83] = 10'b1001101011;
    16'b0110000011010000: out_v[83] = 10'b0110000110;
    16'b0100001011010000: out_v[83] = 10'b1011010110;
    16'b0010001001000000: out_v[83] = 10'b1000011101;
    16'b0000100011010000: out_v[83] = 10'b0001110101;
    16'b0010100011010000: out_v[83] = 10'b1011111001;
    16'b0000000011010000: out_v[83] = 10'b1001111001;
    16'b0000000011000000: out_v[83] = 10'b0100100111;
    16'b0010001011010000: out_v[83] = 10'b1001011001;
    16'b0000001010010000: out_v[83] = 10'b0000100101;
    16'b0010101011010000: out_v[83] = 10'b0100011101;
    16'b0000001011000000: out_v[83] = 10'b1000110001;
    16'b0000001001010000: out_v[83] = 10'b1101000001;
    16'b0000101011010000: out_v[83] = 10'b0110110011;
    16'b0010001011000000: out_v[83] = 10'b1110101001;
    16'b0100000001010000: out_v[83] = 10'b0101000101;
    16'b0000001011100000: out_v[83] = 10'b0001000110;
    16'b0000001001100000: out_v[83] = 10'b0101010101;
    16'b0110100011010000: out_v[83] = 10'b0011001101;
    16'b0010000001010000: out_v[83] = 10'b0111111010;
    16'b0000101010010000: out_v[83] = 10'b1001110011;
    16'b0000000010010000: out_v[83] = 10'b0010011101;
    16'b0010000001100000: out_v[83] = 10'b1111100010;
    16'b0000100010110000: out_v[83] = 10'b0110000110;
    16'b0000000010110000: out_v[83] = 10'b1100011110;
    16'b0000000000100000: out_v[83] = 10'b1100010101;
    16'b0000000000110000: out_v[83] = 10'b1111110100;
    16'b0000000010100000: out_v[83] = 10'b1011100001;
    16'b0110000001100000: out_v[83] = 10'b1001011110;
    16'b0010000000110000: out_v[83] = 10'b0110100010;
    16'b0000000010000000: out_v[83] = 10'b0101110010;
    16'b0110000001110000: out_v[83] = 10'b1000001110;
    16'b0000100010100000: out_v[83] = 10'b1010101010;
    16'b0010000000100000: out_v[83] = 10'b1000111011;
    16'b0010000001110000: out_v[83] = 10'b0010100101;
    16'b0000100000110000: out_v[83] = 10'b1110001010;
    16'b0000000001100000: out_v[83] = 10'b1111010110;
    16'b0100000010110000: out_v[83] = 10'b1001111010;
    16'b0010100000110000: out_v[83] = 10'b0101010111;
    16'b0000000011100000: out_v[83] = 10'b0011010110;
    16'b0010000011110000: out_v[83] = 10'b0101000101;
    16'b0010000011100000: out_v[83] = 10'b0011000111;
    16'b0110000011100000: out_v[83] = 10'b0011110110;
    16'b0010100010110000: out_v[83] = 10'b0101000100;
    16'b0100000011000000: out_v[83] = 10'b1011001110;
    16'b0010000001100001: out_v[83] = 10'b1111100100;
    16'b0100000001100000: out_v[83] = 10'b1100100001;
    16'b0100001001000000: out_v[83] = 10'b1111011001;
    16'b0110001001100000: out_v[83] = 10'b0111011010;
    16'b0110000001010000: out_v[83] = 10'b0111000001;
    16'b0000000001100001: out_v[83] = 10'b1010011110;
    16'b0110000010100000: out_v[83] = 10'b0001101010;
    16'b0100001001100001: out_v[83] = 10'b1110111011;
    16'b0100001011100000: out_v[83] = 10'b1000011110;
    16'b0110001011100000: out_v[83] = 10'b1010110001;
    16'b0100000011100000: out_v[83] = 10'b1001100010;
    16'b0110000011110000: out_v[83] = 10'b0000111011;
    16'b0100000001000000: out_v[83] = 10'b0010110010;
    16'b0100001010100000: out_v[83] = 10'b0001000111;
    16'b0110000011100001: out_v[83] = 10'b1110110110;
    16'b0110001010100000: out_v[83] = 10'b0001100111;
    16'b0100001011000000: out_v[83] = 10'b0100100110;
    16'b0000000011110000: out_v[83] = 10'b0111000100;
    16'b0000000001110000: out_v[83] = 10'b1111010001;
    16'b0100001001100000: out_v[83] = 10'b0110001100;
    16'b0000001010100000: out_v[83] = 10'b1010110110;
    16'b0100000000100000: out_v[83] = 10'b0111000100;
    16'b0010000010100000: out_v[83] = 10'b1100011100;
    16'b0110000011000000: out_v[83] = 10'b0110011111;
    16'b0110001000100000: out_v[83] = 10'b1010000110;
    16'b0110000001100001: out_v[83] = 10'b0111111011;
    16'b0110000001000000: out_v[83] = 10'b1110110101;
    16'b0100001000100000: out_v[83] = 10'b0111001111;
    16'b0010001011100000: out_v[83] = 10'b1010011010;
    16'b0010100011110000: out_v[83] = 10'b0001110111;
    16'b0100000001100001: out_v[83] = 10'b1001000111;
    16'b0100000010100000: out_v[83] = 10'b1101001001;
    16'b0110000000100000: out_v[83] = 10'b0110111101;
    16'b0000100000010000: out_v[83] = 10'b0011100001;
    16'b0000100010010000: out_v[83] = 10'b1001011100;
    16'b0110000010010000: out_v[83] = 10'b1000000111;
    16'b0110001011010000: out_v[83] = 10'b0000011111;
    16'b0100100010010000: out_v[83] = 10'b1001100111;
    16'b0010000000010000: out_v[83] = 10'b1011101010;
    16'b0110100010011000: out_v[83] = 10'b0101110111;
    16'b0000000000010000: out_v[83] = 10'b1000111111;
    16'b0110001011000000: out_v[83] = 10'b1110000101;
    16'b0010100010010000: out_v[83] = 10'b0011001100;
    16'b0110100011110000: out_v[83] = 10'b1010011010;
    16'b0010000001000000: out_v[83] = 10'b1111001010;
    16'b0010000010010000: out_v[83] = 10'b1001110111;
    16'b0000100010011000: out_v[83] = 10'b1100110010;
    16'b0110100010110000: out_v[83] = 10'b0000011111;
    16'b0010001001010000: out_v[83] = 10'b1100011001;
    16'b0110001001010000: out_v[83] = 10'b1010111011;
    16'b0100000010010000: out_v[83] = 10'b0111111000;
    16'b0000000001000001: out_v[83] = 10'b1110110001;
    16'b0110100010010000: out_v[83] = 10'b1111000111;
    16'b0110100010111000: out_v[83] = 10'b0001111110;
    16'b0000100001010000: out_v[83] = 10'b0001001011;
    16'b0110000000000000: out_v[83] = 10'b0000111011;
    16'b0110000000110000: out_v[83] = 10'b0110111011;
    16'b0110000010110000: out_v[83] = 10'b0100110001;
    16'b0010000000000000: out_v[83] = 10'b1111000010;
    16'b0100000000110000: out_v[83] = 10'b0111001011;
    16'b0110100000110000: out_v[83] = 10'b0001111011;
    16'b0110100000000000: out_v[83] = 10'b0101111010;
    16'b0000000000000000: out_v[83] = 10'b0011011110;
    16'b0110000010000000: out_v[83] = 10'b1010000111;
    16'b0100000000010000: out_v[83] = 10'b1111001011;
    16'b0100100000000000: out_v[83] = 10'b1000110100;
    16'b0100000000000000: out_v[83] = 10'b1011010001;
    16'b0110100000100000: out_v[83] = 10'b0011110111;
    16'b0110000000010000: out_v[83] = 10'b0010000010;
    16'b0110100000010000: out_v[83] = 10'b1111000100;
    16'b0100100000010000: out_v[83] = 10'b1101100101;
    16'b0100100010110000: out_v[83] = 10'b0110011001;
    16'b0100100000110000: out_v[83] = 10'b1111000101;
    16'b0100000010000000: out_v[83] = 10'b1111010100;
    16'b0100000010111000: out_v[83] = 10'b1010000011;
    16'b0100100000100000: out_v[83] = 10'b1011101111;
    16'b0100100011110000: out_v[83] = 10'b0110111010;
    16'b0100000001110000: out_v[83] = 10'b1010111001;
    16'b0100000011110000: out_v[83] = 10'b1110001010;
    16'b0110001001000000: out_v[83] = 10'b0010110011;
    16'b0100100010011000: out_v[83] = 10'b1000010100;
    16'b0100100010111000: out_v[83] = 10'b0001101111;
    16'b0100000000100001: out_v[83] = 10'b1011000001;
    16'b0000000000100001: out_v[83] = 10'b0111000000;
    16'b0000000000000001: out_v[83] = 10'b0011100011;
    16'b0010000000100001: out_v[83] = 10'b0100111001;
    16'b0010000010111000: out_v[83] = 10'b0011110111;
    16'b0010100000010000: out_v[83] = 10'b0011000101;
    16'b0000100000011000: out_v[83] = 10'b0011001111;
    16'b0010000000101000: out_v[83] = 10'b0111000101;
    16'b0010100010000000: out_v[83] = 10'b1001000000;
    16'b0000000000111000: out_v[83] = 10'b1000011101;
    16'b0010000010101000: out_v[83] = 10'b0011110101;
    16'b0010100000011000: out_v[83] = 10'b0110001111;
    16'b0000000000011000: out_v[83] = 10'b0110010111;
    16'b0010100010011000: out_v[83] = 10'b1101001000;
    16'b0000000010011000: out_v[83] = 10'b0111001110;
    16'b0010100010000010: out_v[83] = 10'b1101011110;
    16'b0010000010011000: out_v[83] = 10'b1011110011;
    16'b0010000000000010: out_v[83] = 10'b0110101110;
    16'b0010100010010010: out_v[83] = 10'b0111011001;
    16'b0010100000111000: out_v[83] = 10'b0011110110;
    16'b0010000000011000: out_v[83] = 10'b0111100100;
    16'b0010000010000000: out_v[83] = 10'b0110001001;
    16'b0010100010111000: out_v[83] = 10'b1010100011;
    16'b0010000010000010: out_v[83] = 10'b0011110101;
    16'b0010100000000000: out_v[83] = 10'b0000011011;
    16'b0010000011101000: out_v[83] = 10'b0011110001;
    16'b0010100000000010: out_v[83] = 10'b0101001011;
    16'b0000000010101000: out_v[83] = 10'b1100111011;
    16'b0000000010111000: out_v[83] = 10'b1010000001;
    16'b0010000000111000: out_v[83] = 10'b1111010001;
    16'b0010000011111000: out_v[83] = 10'b1001111010;
    16'b0000000000101000: out_v[83] = 10'b1001100110;
    16'b0000000011101000: out_v[83] = 10'b0101111111;
    16'b0010100000010010: out_v[83] = 10'b1011101110;
    16'b0110100011111000: out_v[83] = 10'b0101010000;
    16'b0000100011110000: out_v[83] = 10'b0101010110;
    16'b0010000010110000: out_v[83] = 10'b0011100100;
    16'b0100001011110000: out_v[83] = 10'b0100110110;
    16'b0100100011111000: out_v[83] = 10'b0101110011;
    16'b0000100001110000: out_v[83] = 10'b1101000001;
    16'b0100000000011000: out_v[83] = 10'b1111011010;
    16'b0100000010011000: out_v[83] = 10'b1001101110;
    16'b0010100010100000: out_v[83] = 10'b1111001001;
    16'b0110100010000000: out_v[83] = 10'b1001111101;
    16'b0110100010100000: out_v[83] = 10'b1101101001;
    16'b0000100010111000: out_v[83] = 10'b1111100011;
    16'b0110000000111000: out_v[83] = 10'b1001101110;
    16'b0100000000111000: out_v[83] = 10'b1001100101;
    16'b0110100010000010: out_v[83] = 10'b0111100011;
    16'b0100100010100000: out_v[83] = 10'b1001101001;
    16'b0100000010101000: out_v[83] = 10'b1000100111;
    16'b0110000010000010: out_v[83] = 10'b1100100111;
    16'b0110000010011000: out_v[83] = 10'b0101111111;
    16'b0100100000011000: out_v[83] = 10'b1101100110;
    16'b0110000010100010: out_v[83] = 10'b1101111010;
    16'b0100100010000000: out_v[83] = 10'b0110111101;
    16'b0100000010000010: out_v[83] = 10'b0011101111;
    16'b0110000010111000: out_v[83] = 10'b0011000011;
    default: out_v[83] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010000100001000: out_v[84] = 10'b0100110001;
    16'b0010000100011010: out_v[84] = 10'b0000011011;
    16'b0000000100011000: out_v[84] = 10'b1010101100;
    16'b0010000000001000: out_v[84] = 10'b1101000011;
    16'b0000000101010000: out_v[84] = 10'b1110000011;
    16'b0000000100010000: out_v[84] = 10'b1000001111;
    16'b0000000000011000: out_v[84] = 10'b1111001001;
    16'b0001000001011000: out_v[84] = 10'b1010101111;
    16'b0010000100011000: out_v[84] = 10'b0101010100;
    16'b0010000100001010: out_v[84] = 10'b0011011110;
    16'b0010000000011000: out_v[84] = 10'b1100000110;
    16'b0010000100010010: out_v[84] = 10'b1100100011;
    16'b0010000101011000: out_v[84] = 10'b1110001101;
    16'b0000000101011000: out_v[84] = 10'b1011110110;
    16'b0010000100000000: out_v[84] = 10'b1110100000;
    16'b0010000000001010: out_v[84] = 10'b1110100100;
    16'b0000000000001000: out_v[84] = 10'b1011001110;
    16'b0001000101011000: out_v[84] = 10'b0011011110;
    16'b0000000101001000: out_v[84] = 10'b0011001111;
    16'b0010000001011000: out_v[84] = 10'b1110000111;
    16'b0010000100000010: out_v[84] = 10'b1110110000;
    16'b0010000101011010: out_v[84] = 10'b1110000101;
    16'b0000000100001000: out_v[84] = 10'b0011011010;
    16'b0000000000010000: out_v[84] = 10'b0111011001;
    16'b0000000001011000: out_v[84] = 10'b0001001011;
    16'b0000000100011010: out_v[84] = 10'b1100010011;
    16'b0010000000000000: out_v[84] = 10'b0001011000;
    16'b0000000101011010: out_v[84] = 10'b0110010011;
    16'b0000000001001000: out_v[84] = 10'b0001111111;
    16'b0010000100010000: out_v[84] = 10'b1111001000;
    16'b0000000000000010: out_v[84] = 10'b0110001010;
    16'b0000000100000010: out_v[84] = 10'b1100001101;
    16'b0000000100001010: out_v[84] = 10'b1000111011;
    16'b0000000100000000: out_v[84] = 10'b0010100011;
    16'b0000000000000000: out_v[84] = 10'b0001010010;
    16'b0001000000000010: out_v[84] = 10'b0110001011;
    16'b0010000000000010: out_v[84] = 10'b0001010010;
    16'b0000000000001010: out_v[84] = 10'b1100000000;
    16'b0001000100000000: out_v[84] = 10'b0001110101;
    16'b0001000101001010: out_v[84] = 10'b1011011111;
    16'b0011000001001000: out_v[84] = 10'b1100100011;
    16'b0001000000001000: out_v[84] = 10'b0000110111;
    16'b0001000001001000: out_v[84] = 10'b0010001111;
    16'b0000000101000000: out_v[84] = 10'b1000100100;
    16'b0001000000000000: out_v[84] = 10'b1100010111;
    16'b0001000001000000: out_v[84] = 10'b0011110000;
    16'b0001000101001000: out_v[84] = 10'b1111011011;
    16'b0011000100001000: out_v[84] = 10'b1111000111;
    16'b0011000000001000: out_v[84] = 10'b0110000111;
    16'b0010000101001000: out_v[84] = 10'b0111110011;
    16'b0001000100001010: out_v[84] = 10'b1111011101;
    16'b0011000101001010: out_v[84] = 10'b1001000111;
    16'b0001000100001000: out_v[84] = 10'b1101111100;
    16'b0010000001001000: out_v[84] = 10'b1100101010;
    16'b0010000001001010: out_v[84] = 10'b0110110110;
    16'b0010000101000000: out_v[84] = 10'b1001100110;
    16'b0010000101001010: out_v[84] = 10'b0001101100;
    16'b0000000101001010: out_v[84] = 10'b1101110011;
    16'b0001000101000000: out_v[84] = 10'b1010010110;
    16'b0011000101001000: out_v[84] = 10'b0110010011;
    16'b0000000101000010: out_v[84] = 10'b0101111011;
    16'b0000000001000000: out_v[84] = 10'b1001011111;
    16'b0011000001001010: out_v[84] = 10'b1011100000;
    16'b0011000100001010: out_v[84] = 10'b0010011110;
    16'b0011000000001010: out_v[84] = 10'b1110111110;
    16'b0001000000001010: out_v[84] = 10'b1010100111;
    16'b0010000101000010: out_v[84] = 10'b1110011110;
    16'b0001000100000010: out_v[84] = 10'b0111001000;
    16'b0011000100000010: out_v[84] = 10'b1110100101;
    16'b0010000000010000: out_v[84] = 10'b0001010111;
    16'b0011000000000000: out_v[84] = 10'b1011001001;
    16'b0010000000010010: out_v[84] = 10'b0010101111;
    16'b0010000001000000: out_v[84] = 10'b0101011010;
    16'b0000000001001010: out_v[84] = 10'b0101100000;
    16'b0011000001000000: out_v[84] = 10'b0011000011;
    16'b0001000001010000: out_v[84] = 10'b0111001010;
    16'b0011000000010000: out_v[84] = 10'b1101101111;
    16'b0011000000000010: out_v[84] = 10'b0011001100;
    16'b0001000000010000: out_v[84] = 10'b0111110000;
    16'b0000000001010000: out_v[84] = 10'b0010010011;
    16'b0011000001000010: out_v[84] = 10'b1101101110;
    16'b0010000001000010: out_v[84] = 10'b0011011111;
    16'b0000000010000000: out_v[84] = 10'b1110110011;
    16'b0000000110000000: out_v[84] = 10'b0010110000;
    16'b0000000010000010: out_v[84] = 10'b1110000111;
    16'b0000000110010000: out_v[84] = 10'b1001100111;
    16'b0000000100010010: out_v[84] = 10'b1100110011;
    16'b0000000000010010: out_v[84] = 10'b1011001110;
    16'b0000000000011010: out_v[84] = 10'b1101000110;
    16'b0010000000011010: out_v[84] = 10'b1010001111;
    default: out_v[84] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010000000100000: out_v[85] = 10'b1110010111;
    16'b0010000000110010: out_v[85] = 10'b1010000100;
    16'b0010000000100010: out_v[85] = 10'b0011100101;
    16'b0010000000000010: out_v[85] = 10'b1001101110;
    16'b0000000000100010: out_v[85] = 10'b1101001001;
    16'b0000000000010000: out_v[85] = 10'b0100110101;
    16'b0000000000100000: out_v[85] = 10'b0011110001;
    16'b1010000000100000: out_v[85] = 10'b0111010100;
    16'b0010000010100010: out_v[85] = 10'b0000110111;
    16'b0010000100100010: out_v[85] = 10'b1010100111;
    16'b0010000100110010: out_v[85] = 10'b1011101011;
    16'b0000000100110010: out_v[85] = 10'b1011110011;
    16'b1010000000110010: out_v[85] = 10'b0000010001;
    16'b0000000000110010: out_v[85] = 10'b1100000010;
    16'b0010000000111010: out_v[85] = 10'b0000000101;
    16'b0000000000110000: out_v[85] = 10'b0001011001;
    16'b1010000000100010: out_v[85] = 10'b0010011011;
    16'b0010000110100010: out_v[85] = 10'b0001000111;
    16'b1010000000010010: out_v[85] = 10'b1010001001;
    16'b0010000000010010: out_v[85] = 10'b1000010111;
    16'b0000000000000000: out_v[85] = 10'b0011111001;
    16'b0010000000101010: out_v[85] = 10'b1101010001;
    16'b0000000100100010: out_v[85] = 10'b0010010110;
    16'b0010000010110010: out_v[85] = 10'b1110010011;
    16'b0000000000000010: out_v[85] = 10'b0001111111;
    16'b0010000100000010: out_v[85] = 10'b0001000001;
    16'b0010000000000000: out_v[85] = 10'b0111010011;
    16'b1010000000000010: out_v[85] = 10'b0000011000;
    16'b0010000100000000: out_v[85] = 10'b1011000100;
    16'b1010000000111010: out_v[85] = 10'b1000101111;
    16'b1000000000100000: out_v[85] = 10'b1000000011;
    16'b1000000000101000: out_v[85] = 10'b1001100010;
    16'b1000000000000000: out_v[85] = 10'b1000001010;
    16'b0000000100000000: out_v[85] = 10'b0110011100;
    16'b1000000100000000: out_v[85] = 10'b1000100110;
    16'b1000000110000000: out_v[85] = 10'b1100101011;
    16'b0000000110100000: out_v[85] = 10'b0101100100;
    16'b1000000110100000: out_v[85] = 10'b0110100101;
    16'b0010000100100000: out_v[85] = 10'b1000100110;
    16'b1000000010000000: out_v[85] = 10'b1111000101;
    16'b0000000100100000: out_v[85] = 10'b1000001111;
    16'b0000000110000000: out_v[85] = 10'b1000111100;
    16'b1000000110100001: out_v[85] = 10'b1101100111;
    16'b0000000110000001: out_v[85] = 10'b1011111011;
    16'b1000000100100000: out_v[85] = 10'b0001001001;
    16'b1010000100100000: out_v[85] = 10'b1110001000;
    16'b1010000000000000: out_v[85] = 10'b0110011111;
    16'b0000000000101000: out_v[85] = 10'b0100111110;
    16'b1010000100000000: out_v[85] = 10'b1100010111;
    16'b0000000010000000: out_v[85] = 10'b1001111111;
    16'b0000000000001000: out_v[85] = 10'b0011010001;
    16'b0000000110100001: out_v[85] = 10'b0100011100;
    16'b0000000100100001: out_v[85] = 10'b1110011110;
    16'b0010000110100000: out_v[85] = 10'b1001111100;
    16'b1000000010100000: out_v[85] = 10'b1000011111;
    16'b0000000010100000: out_v[85] = 10'b1000100011;
    16'b1000000110000001: out_v[85] = 10'b0011101101;
    16'b1010000110100000: out_v[85] = 10'b0101000011;
    16'b1010000010000000: out_v[85] = 10'b1110000000;
    16'b0010000010100000: out_v[85] = 10'b0011001000;
    16'b1010000010100000: out_v[85] = 10'b0110011001;
    16'b1010000010100010: out_v[85] = 10'b0010100010;
    16'b1010000010000010: out_v[85] = 10'b1001101010;
    16'b1010000110100010: out_v[85] = 10'b1101001000;
    16'b0010000010000000: out_v[85] = 10'b0010001010;
    16'b1010000110000000: out_v[85] = 10'b1110011010;
    16'b1010000100100010: out_v[85] = 10'b0001011110;
    16'b1000000000000010: out_v[85] = 10'b0010011001;
    16'b0010000010000010: out_v[85] = 10'b0000111100;
    16'b0010000000001000: out_v[85] = 10'b1111011110;
    16'b0000000000010010: out_v[85] = 10'b1110011101;
    16'b0000000010000010: out_v[85] = 10'b0111011011;
    16'b1000000000010000: out_v[85] = 10'b1000100011;
    16'b1010000000101000: out_v[85] = 10'b1101110000;
    16'b0010000000101000: out_v[85] = 10'b1111010010;
    16'b1000000000110000: out_v[85] = 10'b1100100000;
    16'b0000000100000010: out_v[85] = 10'b0111001010;
    16'b1010000100000010: out_v[85] = 10'b0011111010;
    16'b0010000110000010: out_v[85] = 10'b0010010101;
    16'b0010000000001010: out_v[85] = 10'b1011000011;
    16'b0010000100010010: out_v[85] = 10'b0110111010;
    16'b0000100000000000: out_v[85] = 10'b1000001110;
    16'b1000100000000000: out_v[85] = 10'b1111000001;
    16'b0010100000000010: out_v[85] = 10'b0111110010;
    16'b0010100000000000: out_v[85] = 10'b1111000101;
    16'b1010100000000010: out_v[85] = 10'b1011011111;
    default: out_v[85] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010000000000000: out_v[86] = 10'b0001110000;
    16'b0010100000000000: out_v[86] = 10'b0101010001;
    16'b0000000000000000: out_v[86] = 10'b0011001110;
    16'b0000100000000000: out_v[86] = 10'b0000000101;
    16'b0010100000100000: out_v[86] = 10'b0011101011;
    16'b0000000000100000: out_v[86] = 10'b0001011100;
    16'b0010000000100000: out_v[86] = 10'b0110000010;
    16'b0000100000100000: out_v[86] = 10'b1011011011;
    16'b0000000100000000: out_v[86] = 10'b1001000110;
    16'b0000000000001000: out_v[86] = 10'b0011001010;
    16'b0000000000101000: out_v[86] = 10'b0011111101;
    16'b0010000010000000: out_v[86] = 10'b1111100000;
    16'b0010000000001000: out_v[86] = 10'b1001110010;
    16'b0010000100000000: out_v[86] = 10'b0101010111;
    16'b0010000000101000: out_v[86] = 10'b1010011010;
    16'b0010000010100000: out_v[86] = 10'b1111000001;
    16'b0000000010100000: out_v[86] = 10'b1000011110;
    16'b0000000010000000: out_v[86] = 10'b1100101111;
    default: out_v[86] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1000001010100001: out_v[87] = 10'b0101100101;
    16'b0001001010100001: out_v[87] = 10'b0111001011;
    16'b1001001011000001: out_v[87] = 10'b0111111111;
    16'b1000001010000001: out_v[87] = 10'b1110100110;
    16'b0000001010101001: out_v[87] = 10'b1101000000;
    16'b0000001010100001: out_v[87] = 10'b0011100001;
    16'b1001001010101001: out_v[87] = 10'b0111001010;
    16'b1010001010000001: out_v[87] = 10'b1110100001;
    16'b1000001011000000: out_v[87] = 10'b1100011011;
    16'b1011001010000001: out_v[87] = 10'b0010011011;
    16'b0000001000000000: out_v[87] = 10'b1010001011;
    16'b0000000010100001: out_v[87] = 10'b0100111111;
    16'b1011001011000001: out_v[87] = 10'b0001110100;
    16'b1010001011100011: out_v[87] = 10'b0011110101;
    16'b1011001010100001: out_v[87] = 10'b1110010000;
    16'b1000001011000011: out_v[87] = 10'b1011110010;
    16'b1011001011000011: out_v[87] = 10'b0010111011;
    16'b1000001011000001: out_v[87] = 10'b0111011000;
    16'b1010001011000001: out_v[87] = 10'b1101001001;
    16'b1000001000000000: out_v[87] = 10'b1111000010;
    16'b0000001011100001: out_v[87] = 10'b1010111111;
    16'b1000000000000000: out_v[87] = 10'b0100110011;
    16'b1010001011000011: out_v[87] = 10'b0000110010;
    16'b1001001010000001: out_v[87] = 10'b0010010101;
    16'b0001001010101001: out_v[87] = 10'b1000001011;
    16'b0000000000000000: out_v[87] = 10'b0010100101;
    16'b1010001011000010: out_v[87] = 10'b0110101100;
    16'b0000001010000001: out_v[87] = 10'b1100001010;
    16'b0001001000101001: out_v[87] = 10'b0011110001;
    16'b1001001010100001: out_v[87] = 10'b1110001110;
    16'b1000001011100001: out_v[87] = 10'b1011001111;
    16'b0001001010000001: out_v[87] = 10'b0001011101;
    16'b1010001000000000: out_v[87] = 10'b0011011110;
    16'b0000001011000001: out_v[87] = 10'b1110001011;
    16'b1000001010000000: out_v[87] = 10'b1111101010;
    16'b1010001010100001: out_v[87] = 10'b0000110100;
    16'b1010001010000000: out_v[87] = 10'b1001111000;
    16'b1001001011100001: out_v[87] = 10'b1001110111;
    16'b1000001010100000: out_v[87] = 10'b0011110001;
    16'b1000001000100000: out_v[87] = 10'b0011000011;
    16'b0001001011100001: out_v[87] = 10'b1000111110;
    16'b0001001000000000: out_v[87] = 10'b1000001011;
    16'b0001001000001001: out_v[87] = 10'b0001110111;
    16'b0000000010001001: out_v[87] = 10'b0111110100;
    16'b0001001000000001: out_v[87] = 10'b1000001011;
    16'b0000000010000001: out_v[87] = 10'b0100011011;
    16'b0000000000001001: out_v[87] = 10'b0101100111;
    16'b0001001000001000: out_v[87] = 10'b0001010110;
    16'b0001001010001001: out_v[87] = 10'b0010100110;
    16'b0000000000001000: out_v[87] = 10'b0000110111;
    16'b0000001010001001: out_v[87] = 10'b1011101100;
    16'b0001000000000000: out_v[87] = 10'b1100101010;
    16'b0000000010101001: out_v[87] = 10'b0011010001;
    16'b0000001000000001: out_v[87] = 10'b1101011011;
    16'b1000000000001000: out_v[87] = 10'b1001010010;
    16'b0001001000100001: out_v[87] = 10'b1100110011;
    16'b0001000010001001: out_v[87] = 10'b0111101000;
    16'b1000000010001001: out_v[87] = 10'b1101010111;
    16'b1011000010001001: out_v[87] = 10'b0110000100;
    16'b1011001010001101: out_v[87] = 10'b1110011111;
    16'b1011001010001001: out_v[87] = 10'b1000000110;
    16'b1011001000000000: out_v[87] = 10'b0010011110;
    16'b0001000000001000: out_v[87] = 10'b0111101000;
    16'b1001001000001000: out_v[87] = 10'b1100110101;
    16'b1011000000000000: out_v[87] = 10'b1111100100;
    16'b1001001000000000: out_v[87] = 10'b0000110101;
    16'b0010001010001001: out_v[87] = 10'b1101001111;
    16'b1011000000001000: out_v[87] = 10'b0111110110;
    16'b0011001010001001: out_v[87] = 10'b0001011111;
    16'b1010000000001000: out_v[87] = 10'b0001001101;
    16'b1010001010001001: out_v[87] = 10'b1001101100;
    16'b0001001010101011: out_v[87] = 10'b1111101101;
    16'b0001001000101000: out_v[87] = 10'b0001011101;
    16'b1011001010001000: out_v[87] = 10'b0111011001;
    16'b0001001010001011: out_v[87] = 10'b1010001010;
    16'b0010000000001000: out_v[87] = 10'b1000011000;
    16'b1011001010000000: out_v[87] = 10'b1010110011;
    16'b0001001010001000: out_v[87] = 10'b1101100010;
    16'b1011001000001000: out_v[87] = 10'b0111011100;
    16'b0000001010001000: out_v[87] = 10'b1010100010;
    16'b1001001010001001: out_v[87] = 10'b0000111101;
    16'b1000001010001001: out_v[87] = 10'b1101101110;
    16'b0011001000001000: out_v[87] = 10'b0111011011;
    16'b1011001000001100: out_v[87] = 10'b1100111011;
    16'b0000000000101000: out_v[87] = 10'b0100111100;
    16'b1011001010101001: out_v[87] = 10'b0110011101;
    16'b1010001010001000: out_v[87] = 10'b1000001111;
    16'b0000001000001000: out_v[87] = 10'b0111001001;
    16'b1010001000001000: out_v[87] = 10'b0100111010;
    16'b1001001010100000: out_v[87] = 10'b1111000011;
    16'b0001001000100000: out_v[87] = 10'b1100011001;
    16'b0001000000100000: out_v[87] = 10'b0110101001;
    16'b1011001000100000: out_v[87] = 10'b1100000011;
    16'b1001000010100001: out_v[87] = 10'b1001100111;
    16'b1001001000100000: out_v[87] = 10'b0000011000;
    16'b0001001010101000: out_v[87] = 10'b1000001001;
    16'b1001000000100000: out_v[87] = 10'b1110101000;
    16'b1011001010100000: out_v[87] = 10'b0011001100;
    16'b1010000010100001: out_v[87] = 10'b1100011100;
    16'b1011000010100001: out_v[87] = 10'b0010011011;
    16'b0001001010100000: out_v[87] = 10'b1111000111;
    16'b1011000000100000: out_v[87] = 10'b0111011010;
    16'b1010000000100000: out_v[87] = 10'b0000111111;
    16'b1000000010100001: out_v[87] = 10'b0101001100;
    16'b1001001010000000: out_v[87] = 10'b0011111110;
    16'b1000000010000001: out_v[87] = 10'b0100011001;
    16'b0001001010000000: out_v[87] = 10'b0011011111;
    16'b1001001000100001: out_v[87] = 10'b0101011110;
    16'b1011001000100001: out_v[87] = 10'b0110011101;
    16'b0001000000101000: out_v[87] = 10'b0010111101;
    16'b1001001010101000: out_v[87] = 10'b1110001111;
    16'b1001001000101000: out_v[87] = 10'b0110010010;
    16'b0000000000101001: out_v[87] = 10'b1000101111;
    16'b1000000000100000: out_v[87] = 10'b1010100111;
    16'b1001000000101000: out_v[87] = 10'b0101000000;
    16'b0000000000100000: out_v[87] = 10'b0101111011;
    16'b1000000000101000: out_v[87] = 10'b1110011111;
    16'b1001000000001000: out_v[87] = 10'b1011101011;
    16'b0001000010101001: out_v[87] = 10'b1001110100;
    16'b0001000000101001: out_v[87] = 10'b1010001000;
    16'b1011001000101000: out_v[87] = 10'b1010000111;
    16'b1010001010100000: out_v[87] = 10'b1010100011;
    16'b0000001000101001: out_v[87] = 10'b0100101011;
    16'b1000001010101001: out_v[87] = 10'b1011100101;
    16'b1000000010100000: out_v[87] = 10'b0110110011;
    16'b0000001010100000: out_v[87] = 10'b0101100110;
    16'b0001000000100001: out_v[87] = 10'b0111111000;
    16'b1010000010100000: out_v[87] = 10'b0010100001;
    16'b0000001000100001: out_v[87] = 10'b1001011001;
    16'b1010001010101001: out_v[87] = 10'b0011100110;
    16'b0000000010100000: out_v[87] = 10'b0111111000;
    16'b0000100000000000: out_v[87] = 10'b1111110111;
    16'b1000000010101000: out_v[87] = 10'b0011001101;
    16'b1000100000100000: out_v[87] = 10'b1111001100;
    16'b1000000010101001: out_v[87] = 10'b0100010111;
    16'b0000100000101000: out_v[87] = 10'b1101110011;
    16'b1000100000101000: out_v[87] = 10'b0011101101;
    16'b1000100000001000: out_v[87] = 10'b1110111001;
    16'b0000100000001000: out_v[87] = 10'b0000111111;
    16'b0000000010101000: out_v[87] = 10'b0100111010;
    16'b1010000000000000: out_v[87] = 10'b0111110110;
    16'b0000100000100000: out_v[87] = 10'b1011011010;
    16'b0000000000001100: out_v[87] = 10'b0110100001;
    16'b0001000000001001: out_v[87] = 10'b1110000000;
    16'b1001000000000000: out_v[87] = 10'b0110101000;
    16'b1001000000001001: out_v[87] = 10'b1001111011;
    16'b0001000000000001: out_v[87] = 10'b1011100000;
    16'b1001000000000001: out_v[87] = 10'b0011100110;
    16'b0000001000001001: out_v[87] = 10'b1111000001;
    16'b1000001010101000: out_v[87] = 10'b1110100011;
    16'b0000001010101000: out_v[87] = 10'b1111100010;
    16'b0001000010101000: out_v[87] = 10'b1000011010;
    16'b1001000010101001: out_v[87] = 10'b1001100010;
    16'b1001000010000001: out_v[87] = 10'b1000000101;
    16'b0001000010000001: out_v[87] = 10'b0101001101;
    16'b1001000010001001: out_v[87] = 10'b1000101001;
    default: out_v[87] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010001000100011: out_v[88] = 10'b0010111111;
    16'b0000001000101111: out_v[88] = 10'b1110011110;
    16'b0010101100101111: out_v[88] = 10'b0100001101;
    16'b0010101000101011: out_v[88] = 10'b0010100110;
    16'b0000001000101011: out_v[88] = 10'b0010100111;
    16'b0000100100101011: out_v[88] = 10'b1000110010;
    16'b0010001000111101: out_v[88] = 10'b1011111010;
    16'b0010001000101001: out_v[88] = 10'b1000110011;
    16'b0010001000101101: out_v[88] = 10'b1110101111;
    16'b0000001000111111: out_v[88] = 10'b0001111000;
    16'b0010001000101011: out_v[88] = 10'b1110100011;
    16'b0010100000101011: out_v[88] = 10'b0000111011;
    16'b0010101100101011: out_v[88] = 10'b1010111001;
    16'b0010001000101111: out_v[88] = 10'b1110011011;
    16'b0010101100111101: out_v[88] = 10'b0001000101;
    16'b0010101000101111: out_v[88] = 10'b0110011011;
    16'b0010101100100010: out_v[88] = 10'b1011111101;
    16'b0000000000101111: out_v[88] = 10'b1100001010;
    16'b0010101000100010: out_v[88] = 10'b1010111110;
    16'b0000001000111101: out_v[88] = 10'b1100110110;
    16'b0010101100101101: out_v[88] = 10'b0101010000;
    16'b0000000000111101: out_v[88] = 10'b0010011010;
    16'b0000101000101011: out_v[88] = 10'b1010000101;
    16'b0010101100111111: out_v[88] = 10'b1111100111;
    16'b0010101100101010: out_v[88] = 10'b0010110011;
    16'b0010001100101011: out_v[88] = 10'b1100011011;
    16'b0010001000001011: out_v[88] = 10'b1000011011;
    16'b0010100100101011: out_v[88] = 10'b0111100111;
    16'b0010101000101001: out_v[88] = 10'b0010110110;
    16'b0010001100101111: out_v[88] = 10'b0111101110;
    16'b0010001100111101: out_v[88] = 10'b1111111111;
    16'b0010100000100010: out_v[88] = 10'b1111110111;
    16'b0010001000111111: out_v[88] = 10'b1011001011;
    16'b0000001010100000: out_v[88] = 10'b1001101111;
    16'b0010000010001000: out_v[88] = 10'b0101110110;
    16'b0010000010001001: out_v[88] = 10'b0011100111;
    16'b0000001010000000: out_v[88] = 10'b1000001100;
    16'b0010000010000000: out_v[88] = 10'b0011011011;
    16'b0010000010000001: out_v[88] = 10'b0100110000;
    16'b0000000010100000: out_v[88] = 10'b1001010111;
    16'b0000001010001000: out_v[88] = 10'b0100111111;
    16'b0010001010100000: out_v[88] = 10'b1101001101;
    16'b0000000010000000: out_v[88] = 10'b1011000100;
    16'b0000000010001001: out_v[88] = 10'b0011011110;
    16'b0000100010000001: out_v[88] = 10'b0111110011;
    16'b0010001010001000: out_v[88] = 10'b1111001000;
    16'b0000000010000001: out_v[88] = 10'b1101001001;
    16'b0000001010101000: out_v[88] = 10'b0010001010;
    16'b0000100010001001: out_v[88] = 10'b0010110011;
    16'b0000001000000000: out_v[88] = 10'b1010110010;
    16'b0010001010101000: out_v[88] = 10'b0110101011;
    16'b0010001010001001: out_v[88] = 10'b1111011110;
    16'b0010000000001000: out_v[88] = 10'b0111010010;
    16'b0000000010001000: out_v[88] = 10'b1010010100;
    16'b0000000010100100: out_v[88] = 10'b1011011111;
    16'b0010100010001001: out_v[88] = 10'b1101001011;
    16'b0000001010001001: out_v[88] = 10'b1001010100;
    16'b0000001010101001: out_v[88] = 10'b1011000010;
    16'b0010001010101001: out_v[88] = 10'b0011111100;
    16'b0010100010101001: out_v[88] = 10'b0101011011;
    16'b0010000010101001: out_v[88] = 10'b1111011001;
    16'b0010101010101001: out_v[88] = 10'b0000111010;
    16'b0000101010101001: out_v[88] = 10'b1100100111;
    16'b0000101010100000: out_v[88] = 10'b0100000111;
    16'b0010100010000000: out_v[88] = 10'b0011101000;
    16'b0010101010100001: out_v[88] = 10'b1011010011;
    16'b0010101010100011: out_v[88] = 10'b0101011110;
    16'b0000001000101001: out_v[88] = 10'b0011001000;
    16'b0000001010000001: out_v[88] = 10'b0100010101;
    16'b0010101010100010: out_v[88] = 10'b1110000101;
    16'b0010101010100000: out_v[88] = 10'b0001010100;
    16'b0010001010100001: out_v[88] = 10'b0100100100;
    16'b0010101010000001: out_v[88] = 10'b1011101000;
    16'b0010100000101001: out_v[88] = 10'b1100011100;
    16'b0000101000101001: out_v[88] = 10'b0111110010;
    16'b0010100010100001: out_v[88] = 10'b1110000101;
    16'b0000101010100001: out_v[88] = 10'b1010001011;
    16'b0010101010101011: out_v[88] = 10'b0000011110;
    16'b0010000000101001: out_v[88] = 10'b0001011011;
    16'b0010101000100011: out_v[88] = 10'b0101001010;
    16'b0000001010100001: out_v[88] = 10'b1111001000;
    16'b0010001010100111: out_v[88] = 10'b1011111111;
    16'b0010001010100010: out_v[88] = 10'b1011100110;
    16'b0010001010101011: out_v[88] = 10'b0011000011;
    16'b0010101010101111: out_v[88] = 10'b1001111110;
    16'b0010101010101000: out_v[88] = 10'b0010111011;
    16'b0010001010000001: out_v[88] = 10'b1101001001;
    16'b0000100010000000: out_v[88] = 10'b1000001100;
    16'b0010100010000001: out_v[88] = 10'b1100000101;
    16'b0010100010100000: out_v[88] = 10'b0110110000;
    16'b0010001010000000: out_v[88] = 10'b1110000001;
    16'b0010000010100000: out_v[88] = 10'b0010111111;
    16'b0010101010001001: out_v[88] = 10'b1001101001;
    16'b0010101010000000: out_v[88] = 10'b1110011000;
    16'b0010001010101111: out_v[88] = 10'b1010010110;
    16'b0000100010101001: out_v[88] = 10'b0011100110;
    16'b0010101000001001: out_v[88] = 10'b0111101110;
    16'b0010101010001111: out_v[88] = 10'b0101011011;
    16'b0000101010000001: out_v[88] = 10'b0111010100;
    16'b0000000010001110: out_v[88] = 10'b1000101011;
    16'b0000100010001000: out_v[88] = 10'b0110111001;
    16'b0000100010000011: out_v[88] = 10'b1101101001;
    16'b0000000110000001: out_v[88] = 10'b0111011011;
    16'b0000000010000110: out_v[88] = 10'b1011001110;
    16'b0100000110000000: out_v[88] = 10'b1100111111;
    16'b0000000010100110: out_v[88] = 10'b1000011011;
    16'b0000100110000011: out_v[88] = 10'b0101101010;
    16'b0000100010001011: out_v[88] = 10'b1101111111;
    16'b0000100110001001: out_v[88] = 10'b0011110110;
    16'b0000100000000011: out_v[88] = 10'b0011011111;
    16'b0000101000000001: out_v[88] = 10'b0001111010;
    16'b0000001110000001: out_v[88] = 10'b0001011011;
    16'b0000101010001001: out_v[88] = 10'b0001011011;
    16'b0000100000000001: out_v[88] = 10'b0111000110;
    16'b0000000000000001: out_v[88] = 10'b0100111110;
    16'b0000100010001111: out_v[88] = 10'b0011011011;
    16'b0000000010001111: out_v[88] = 10'b1101001110;
    16'b0000100110001011: out_v[88] = 10'b0011111111;
    16'b0000100110001111: out_v[88] = 10'b0110011111;
    16'b0000001000000001: out_v[88] = 10'b0111011101;
    16'b0000100110000001: out_v[88] = 10'b1100101110;
    16'b0000000110001001: out_v[88] = 10'b1001110100;
    16'b0000000010111101: out_v[88] = 10'b0000100111;
    16'b0010101010101101: out_v[88] = 10'b1000110111;
    16'b0000000000101101: out_v[88] = 10'b1110110110;
    16'b0000000010101101: out_v[88] = 10'b1110000111;
    16'b0000000010110100: out_v[88] = 10'b1101111000;
    16'b0000000010010100: out_v[88] = 10'b0111100000;
    16'b0000000010101001: out_v[88] = 10'b0110101100;
    16'b0010001010101101: out_v[88] = 10'b1011100110;
    16'b0010101000000000: out_v[88] = 10'b1000100111;
    16'b0010001000001001: out_v[88] = 10'b1011100101;
    16'b0000000010001101: out_v[88] = 10'b1011100111;
    16'b0010101000100000: out_v[88] = 10'b1000011011;
    16'b0000000000100100: out_v[88] = 10'b1011111100;
    16'b0000000010000100: out_v[88] = 10'b0010110000;
    16'b0000100010101101: out_v[88] = 10'b1101010111;
    16'b0000000000110100: out_v[88] = 10'b1001010101;
    16'b0010101000100001: out_v[88] = 10'b1101011001;
    16'b0000000000101001: out_v[88] = 10'b0111110100;
    16'b0010101110101001: out_v[88] = 10'b0000110110;
    16'b0000100010101011: out_v[88] = 10'b0011000001;
    16'b0000100000001001: out_v[88] = 10'b0001011010;
    16'b0010000000001001: out_v[88] = 10'b1011000010;
    16'b0000100110101011: out_v[88] = 10'b1101100010;
    16'b0010000010101011: out_v[88] = 10'b0101000000;
    16'b0010100010101011: out_v[88] = 10'b1100101110;
    16'b0000001000001001: out_v[88] = 10'b0110110011;
    16'b0000000000001001: out_v[88] = 10'b0011110100;
    16'b0000100000001011: out_v[88] = 10'b0011001010;
    16'b0000000100000011: out_v[88] = 10'b0011101011;
    16'b0000100010100010: out_v[88] = 10'b0011110111;
    16'b0000000110001000: out_v[88] = 10'b0110001100;
    16'b0000000100001001: out_v[88] = 10'b0001011110;
    16'b0000100010001010: out_v[88] = 10'b0101110111;
    16'b0000000100001111: out_v[88] = 10'b1101011110;
    16'b0000100010100000: out_v[88] = 10'b0010010000;
    16'b0010100010001000: out_v[88] = 10'b1110000000;
    16'b0000000010001010: out_v[88] = 10'b1100001010;
    16'b0000100100001011: out_v[88] = 10'b0101011101;
    16'b0000000000001000: out_v[88] = 10'b1001101110;
    16'b0000000100000010: out_v[88] = 10'b1100000001;
    16'b0000000010100010: out_v[88] = 10'b1010000110;
    16'b0000000000001010: out_v[88] = 10'b0011111010;
    16'b0000000000001011: out_v[88] = 10'b0111000010;
    16'b0000000100000001: out_v[88] = 10'b1110001011;
    16'b0000100000001010: out_v[88] = 10'b1010101011;
    16'b0000100100001111: out_v[88] = 10'b0011111001;
    16'b0000000000000011: out_v[88] = 10'b1010001111;
    16'b0000000100001011: out_v[88] = 10'b0111000000;
    16'b0000100100000011: out_v[88] = 10'b0100011111;
    16'b0000100010100110: out_v[88] = 10'b1001011011;
    16'b0000000110001011: out_v[88] = 10'b1001100110;
    16'b0010001010111111: out_v[88] = 10'b0111001000;
    16'b0000000010110110: out_v[88] = 10'b1101000110;
    16'b0010101010111111: out_v[88] = 10'b1011111101;
    16'b0010101010100111: out_v[88] = 10'b1010101011;
    16'b0010101010011111: out_v[88] = 10'b1010101110;
    16'b0010001010001111: out_v[88] = 10'b1011011111;
    16'b0010100010001011: out_v[88] = 10'b1001111011;
    16'b0010100110000011: out_v[88] = 10'b1001101000;
    16'b0110100110000000: out_v[88] = 10'b1010100011;
    16'b0000000010001011: out_v[88] = 10'b1011101011;
    16'b0010100000000001: out_v[88] = 10'b1011001011;
    16'b0110100110000010: out_v[88] = 10'b1010100011;
    16'b0110100110000001: out_v[88] = 10'b1111100111;
    16'b0000000010000010: out_v[88] = 10'b1011101100;
    16'b0100100110000000: out_v[88] = 10'b0001011001;
    16'b0010000010001011: out_v[88] = 10'b0110111001;
    16'b0010100110000001: out_v[88] = 10'b1011010111;
    16'b0010100110001011: out_v[88] = 10'b1101001111;
    16'b0010000010001010: out_v[88] = 10'b1011001011;
    16'b0000000110000011: out_v[88] = 10'b1001010001;
    default: out_v[88] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000001000000000: out_v[89] = 10'b0111110010;
    16'b0000101000000000: out_v[89] = 10'b0011100011;
    16'b0001101000000000: out_v[89] = 10'b0101011001;
    16'b0001001000000000: out_v[89] = 10'b1010100110;
    16'b0010001000000000: out_v[89] = 10'b0101010001;
    16'b0101101000000000: out_v[89] = 10'b0111011111;
    16'b0010100000010000: out_v[89] = 10'b1011010001;
    16'b0010101000010000: out_v[89] = 10'b1101011110;
    16'b1101100000000000: out_v[89] = 10'b0101100100;
    16'b0010101000000000: out_v[89] = 10'b0111010100;
    16'b0000100000000000: out_v[89] = 10'b1010100011;
    16'b1001000000000000: out_v[89] = 10'b0110100011;
    16'b0001100000000000: out_v[89] = 10'b1100010111;
    16'b0010000000010000: out_v[89] = 10'b1001111010;
    16'b1101101000000000: out_v[89] = 10'b0110000101;
    16'b1001100000000000: out_v[89] = 10'b1111010111;
    16'b1001101000000000: out_v[89] = 10'b1001010100;
    16'b0101100000000000: out_v[89] = 10'b0100011010;
    16'b0001000000000000: out_v[89] = 10'b1000011001;
    16'b0111101000010000: out_v[89] = 10'b0010100111;
    16'b0010000000000000: out_v[89] = 10'b0101010011;
    16'b0010001000010000: out_v[89] = 10'b0101111000;
    16'b0100101000000000: out_v[89] = 10'b1000010001;
    16'b0011101000000000: out_v[89] = 10'b0010010011;
    16'b0100100000000000: out_v[89] = 10'b1000001011;
    16'b0000000000000000: out_v[89] = 10'b0011100111;
    16'b1001001000000000: out_v[89] = 10'b0010100001;
    16'b0011101000010000: out_v[89] = 10'b1110011100;
    16'b0101000000000000: out_v[89] = 10'b0101001011;
    16'b0000000000010000: out_v[89] = 10'b1110010010;
    16'b1010000000010000: out_v[89] = 10'b1110110100;
    16'b0011000000010000: out_v[89] = 10'b0111011000;
    16'b1010000000000000: out_v[89] = 10'b0100001011;
    16'b1011000000010000: out_v[89] = 10'b1111100100;
    16'b1011001000010000: out_v[89] = 10'b1001100110;
    16'b1111001000010000: out_v[89] = 10'b0101011000;
    16'b1000001000000000: out_v[89] = 10'b1010001000;
    16'b0111001010010000: out_v[89] = 10'b0010010110;
    16'b1010010000010000: out_v[89] = 10'b0011111000;
    16'b0110000000010000: out_v[89] = 10'b0110110000;
    16'b1111000010010000: out_v[89] = 10'b0111110011;
    16'b1000000000000000: out_v[89] = 10'b0000001001;
    16'b0011001000010000: out_v[89] = 10'b0100011001;
    16'b0111001000010000: out_v[89] = 10'b0001010110;
    16'b0110001000010000: out_v[89] = 10'b0001010100;
    16'b1111001010010000: out_v[89] = 10'b0111000100;
    16'b1010011000010000: out_v[89] = 10'b1100110000;
    16'b0111000010010000: out_v[89] = 10'b1000000100;
    16'b1011001010010000: out_v[89] = 10'b0011001110;
    16'b1110000000010000: out_v[89] = 10'b1110100011;
    16'b1111011000010000: out_v[89] = 10'b1110110101;
    16'b1010001000010000: out_v[89] = 10'b1000101011;
    16'b0011100000010000: out_v[89] = 10'b1110010100;
    16'b0011001010010000: out_v[89] = 10'b0100110100;
    16'b0111000000010000: out_v[89] = 10'b1001010110;
    16'b1110011000010000: out_v[89] = 10'b1010110101;
    16'b1111000000010000: out_v[89] = 10'b0011010100;
    16'b0001000000010000: out_v[89] = 10'b1100100100;
    16'b1011101000010000: out_v[89] = 10'b0011110001;
    16'b1001000000010000: out_v[89] = 10'b1101010110;
    16'b0001001000100000: out_v[89] = 10'b1101010100;
    16'b0001000000100000: out_v[89] = 10'b0000101000;
    16'b1010001000000000: out_v[89] = 10'b0011001110;
    16'b0011001000000000: out_v[89] = 10'b1001001000;
    16'b0011000000000000: out_v[89] = 10'b1011001010;
    16'b0001001000000001: out_v[89] = 10'b0100011111;
    16'b1100000000000000: out_v[89] = 10'b0001101011;
    16'b1101000000000000: out_v[89] = 10'b1010101110;
    16'b0010000100010000: out_v[89] = 10'b1011110000;
    16'b0011000000100000: out_v[89] = 10'b1110100000;
    16'b0000000000100000: out_v[89] = 10'b1101010111;
    16'b0010000000100000: out_v[89] = 10'b1111101001;
    16'b0001000100000000: out_v[89] = 10'b1010110100;
    16'b0001001100000000: out_v[89] = 10'b1100000011;
    16'b0000001100000000: out_v[89] = 10'b0100110110;
    16'b0010000100000000: out_v[89] = 10'b1111111010;
    16'b1111111000010000: out_v[89] = 10'b0111111111;
    16'b1011111000010000: out_v[89] = 10'b0100001110;
    16'b0000001000010000: out_v[89] = 10'b0111000101;
    16'b1111101000010000: out_v[89] = 10'b1001100010;
    16'b1011011000010000: out_v[89] = 10'b1010001001;
    16'b0000001000100000: out_v[89] = 10'b1101000011;
    16'b0011001000100000: out_v[89] = 10'b1101110011;
    16'b0011001000110000: out_v[89] = 10'b0100111000;
    16'b0011000000110000: out_v[89] = 10'b0010010101;
    16'b0010000000110000: out_v[89] = 10'b0110111011;
    16'b0000001000001000: out_v[89] = 10'b0011000011;
    16'b0010001000100000: out_v[89] = 10'b0101101110;
    16'b0000101000100000: out_v[89] = 10'b0011011110;
    16'b0000001000101000: out_v[89] = 10'b0111011110;
    16'b0001001000010000: out_v[89] = 10'b1000110111;
    16'b0010100000000000: out_v[89] = 10'b1100011011;
    16'b0010001000110000: out_v[89] = 10'b1001001010;
    default: out_v[89] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1010000000011000: out_v[90] = 10'b1011010101;
    16'b1010000000001000: out_v[90] = 10'b1001101010;
    16'b1010010000001000: out_v[90] = 10'b1001000001;
    16'b1000010000001000: out_v[90] = 10'b0010100011;
    16'b1000010000001010: out_v[90] = 10'b1010011001;
    16'b1010000000010000: out_v[90] = 10'b0110111100;
    16'b1000010000000000: out_v[90] = 10'b0001011011;
    16'b1010010000001010: out_v[90] = 10'b0001010111;
    16'b0000010000001010: out_v[90] = 10'b1000000111;
    16'b1010000000000000: out_v[90] = 10'b1100101111;
    16'b0010010000001000: out_v[90] = 10'b0101110010;
    16'b0010000000011000: out_v[90] = 10'b0001011011;
    16'b1010010000011000: out_v[90] = 10'b0101000001;
    16'b1000010000000010: out_v[90] = 10'b1001101111;
    16'b0010000000001000: out_v[90] = 10'b0011110111;
    16'b1000000000011000: out_v[90] = 10'b0100101010;
    16'b1010010000010000: out_v[90] = 10'b1100110010;
    16'b1000000000000000: out_v[90] = 10'b0000111001;
    16'b0000010000000000: out_v[90] = 10'b0111000010;
    16'b1000010000011000: out_v[90] = 10'b0110100100;
    16'b1000000000010000: out_v[90] = 10'b0101010001;
    16'b1010010000000000: out_v[90] = 10'b1000101000;
    16'b0010000000000000: out_v[90] = 10'b1001101011;
    16'b0010010000001010: out_v[90] = 10'b0011010111;
    16'b0000010000001000: out_v[90] = 10'b1000010100;
    16'b1000000000001000: out_v[90] = 10'b0100110000;
    16'b0000000000000000: out_v[90] = 10'b1101001010;
    16'b0000000010000000: out_v[90] = 10'b1010000001;
    16'b0000000000001000: out_v[90] = 10'b1000001110;
    16'b0000000000011000: out_v[90] = 10'b1010011100;
    16'b0010000000010000: out_v[90] = 10'b0110111100;
    16'b0000000000010000: out_v[90] = 10'b1011110010;
    16'b0010010000011000: out_v[90] = 10'b0111001011;
    16'b0000010000010000: out_v[90] = 10'b0111111011;
    16'b0010000000011010: out_v[90] = 10'b1001011010;
    16'b1000010000010000: out_v[90] = 10'b0100001011;
    16'b0000010000011000: out_v[90] = 10'b1100010110;
    16'b0000000000011010: out_v[90] = 10'b0001101110;
    16'b0000000000001010: out_v[90] = 10'b0101100001;
    16'b0000010000011010: out_v[90] = 10'b0111100011;
    16'b0010000000001010: out_v[90] = 10'b0111000111;
    16'b0010010000010000: out_v[90] = 10'b1101010001;
    16'b1000010000010100: out_v[90] = 10'b0011001101;
    16'b1000000001010000: out_v[90] = 10'b0111110101;
    16'b1000000010000000: out_v[90] = 10'b0001011011;
    16'b1000000010010000: out_v[90] = 10'b0100100011;
    16'b1000010010010000: out_v[90] = 10'b1010111110;
    16'b0010010000011010: out_v[90] = 10'b0011110001;
    16'b0010010000000000: out_v[90] = 10'b1001100010;
    16'b0010000000010100: out_v[90] = 10'b0001110111;
    16'b0000010000010100: out_v[90] = 10'b0010000111;
    16'b0000010010010000: out_v[90] = 10'b0010001011;
    16'b0000010000000100: out_v[90] = 10'b0011011101;
    16'b0000000010010000: out_v[90] = 10'b0011000011;
    default: out_v[90] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000100001100000: out_v[91] = 10'b0110000011;
    16'b0000100001100010: out_v[91] = 10'b1001100001;
    16'b0000110001101010: out_v[91] = 10'b1000000101;
    16'b0000110000101010: out_v[91] = 10'b1100001010;
    16'b0000100000100000: out_v[91] = 10'b0111101011;
    16'b0000010001001000: out_v[91] = 10'b0110011001;
    16'b0000110000001010: out_v[91] = 10'b1000001001;
    16'b0000110000000000: out_v[91] = 10'b1010011111;
    16'b0000100000000000: out_v[91] = 10'b0111010011;
    16'b0000110001101000: out_v[91] = 10'b0011000111;
    16'b0000110000100010: out_v[91] = 10'b1110101010;
    16'b0000110001100010: out_v[91] = 10'b0010111101;
    16'b0000010000101000: out_v[91] = 10'b0110110000;
    16'b0000100001101000: out_v[91] = 10'b1100000100;
    16'b0000000001100000: out_v[91] = 10'b1011001001;
    16'b0000100000100010: out_v[91] = 10'b1101000111;
    16'b0000110000101000: out_v[91] = 10'b0001110010;
    16'b0000110001001000: out_v[91] = 10'b1001110000;
    16'b0000010001100000: out_v[91] = 10'b0111011111;
    16'b0000110001001010: out_v[91] = 10'b0100010111;
    16'b0000010000001000: out_v[91] = 10'b0011001010;
    16'b0000100001000000: out_v[91] = 10'b1100100000;
    16'b0000100001000010: out_v[91] = 10'b0100110100;
    16'b0000010000101010: out_v[91] = 10'b0001100001;
    16'b0000110000001000: out_v[91] = 10'b0000111011;
    16'b1000110001101000: out_v[91] = 10'b0011110011;
    16'b0000100001101010: out_v[91] = 10'b1100111011;
    16'b0000100000101000: out_v[91] = 10'b0101011010;
    16'b0000000000100000: out_v[91] = 10'b0010110111;
    16'b0000100000101010: out_v[91] = 10'b0111101001;
    16'b0000000000000000: out_v[91] = 10'b1100100000;
    16'b1000100001100010: out_v[91] = 10'b1110101101;
    16'b1000100001100000: out_v[91] = 10'b0011101011;
    16'b0000000001000000: out_v[91] = 10'b1111001101;
    16'b0000110001100000: out_v[91] = 10'b0110011011;
    16'b0000110000100000: out_v[91] = 10'b1110001001;
    16'b0000010001101000: out_v[91] = 10'b1010010011;
    16'b0000010000100000: out_v[91] = 10'b0011100100;
    16'b1000100001101000: out_v[91] = 10'b1000111110;
    16'b1000100001101010: out_v[91] = 10'b1101000011;
    16'b1000110001101010: out_v[91] = 10'b0011011110;
    16'b1000100000000010: out_v[91] = 10'b1001100111;
    16'b1000100000000000: out_v[91] = 10'b0111110000;
    16'b1000000001000000: out_v[91] = 10'b0011010010;
    16'b1000000000000000: out_v[91] = 10'b1100010101;
    16'b0000100000000010: out_v[91] = 10'b0010001010;
    16'b1000000000000010: out_v[91] = 10'b1100011000;
    16'b1000100001000000: out_v[91] = 10'b0111000100;
    16'b1000100001000010: out_v[91] = 10'b1001100110;
    16'b1000100000001000: out_v[91] = 10'b0101011000;
    16'b1000000000010000: out_v[91] = 10'b1101111111;
    16'b1000100000100000: out_v[91] = 10'b1101001111;
    16'b1000110000100000: out_v[91] = 10'b0100110110;
    16'b1000100000101000: out_v[91] = 10'b1000011011;
    16'b1000010000100000: out_v[91] = 10'b1111100100;
    16'b1000000000100000: out_v[91] = 10'b0001000001;
    16'b1000110000000000: out_v[91] = 10'b0110110110;
    16'b1000100000100010: out_v[91] = 10'b0010011001;
    16'b1000010000000000: out_v[91] = 10'b0111110011;
    16'b1000010001000000: out_v[91] = 10'b1100110110;
    16'b1000010001010000: out_v[91] = 10'b1100110101;
    16'b1000010001110000: out_v[91] = 10'b1110001110;
    16'b1000010001100000: out_v[91] = 10'b0110101111;
    16'b0000000000000010: out_v[91] = 10'b0101110000;
    16'b1000110000100010: out_v[91] = 10'b0110111010;
    16'b1000000001010000: out_v[91] = 10'b1110101110;
    16'b0000000000100010: out_v[91] = 10'b0111110001;
    16'b0000000001000010: out_v[91] = 10'b0110001000;
    16'b0000010001100010: out_v[91] = 10'b1011011110;
    16'b0000010000100010: out_v[91] = 10'b0110100001;
    16'b0000000001100010: out_v[91] = 10'b0111011011;
    16'b0000000000001000: out_v[91] = 10'b0111110011;
    16'b0000000000101000: out_v[91] = 10'b1010001100;
    16'b1000110000101000: out_v[91] = 10'b1000111011;
    16'b0000100000001000: out_v[91] = 10'b1011101010;
    16'b1000000000001000: out_v[91] = 10'b0111001100;
    16'b1000000000101000: out_v[91] = 10'b0001011000;
    16'b1000000001000010: out_v[91] = 10'b0010010110;
    16'b1000010000101000: out_v[91] = 10'b0101010001;
    16'b0000000001101000: out_v[91] = 10'b1110100110;
    16'b0000100001001010: out_v[91] = 10'b1000100011;
    16'b0000100001001000: out_v[91] = 10'b0010100011;
    16'b0000000001001000: out_v[91] = 10'b1111100001;
    16'b1000000001100000: out_v[91] = 10'b1111101010;
    16'b1000010000111000: out_v[91] = 10'b0011001011;
    16'b1000000000000100: out_v[91] = 10'b1100011001;
    16'b1000010000100100: out_v[91] = 10'b1010011101;
    16'b1000010000001000: out_v[91] = 10'b0001000011;
    16'b0000000000100100: out_v[91] = 10'b1111111110;
    16'b0000010000100100: out_v[91] = 10'b1100110110;
    16'b1000000000100100: out_v[91] = 10'b1110100101;
    16'b0000010000000000: out_v[91] = 10'b1011100010;
    16'b1000010000101100: out_v[91] = 10'b1000110011;
    16'b1000010001101000: out_v[91] = 10'b1110000011;
    16'b1000100001001000: out_v[91] = 10'b1101010110;
    16'b1000000001100010: out_v[91] = 10'b0010011100;
    16'b1000000001101000: out_v[91] = 10'b1100100111;
    default: out_v[91] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1001110000000000: out_v[92] = 10'b0110011111;
    16'b0001100010010001: out_v[92] = 10'b1111111111;
    16'b0001110010010000: out_v[92] = 10'b0101111111;
    16'b1001100010000001: out_v[92] = 10'b1000101111;
    16'b1001110010000001: out_v[92] = 10'b0010100111;
    16'b1001110010010000: out_v[92] = 10'b0000001101;
    16'b1001110011010000: out_v[92] = 10'b0011000111;
    16'b0000000000000001: out_v[92] = 10'b0001110011;
    16'b1001111000010000: out_v[92] = 10'b0010001001;
    16'b0000110010000001: out_v[92] = 10'b1010011101;
    16'b1001110010010001: out_v[92] = 10'b0010010100;
    16'b0000100010000001: out_v[92] = 10'b1000010111;
    16'b1001100010010000: out_v[92] = 10'b0111110111;
    16'b0000000010000001: out_v[92] = 10'b1101011110;
    16'b0001110010000000: out_v[92] = 10'b0100010111;
    16'b1001111010010000: out_v[92] = 10'b1001000111;
    16'b0000100010000000: out_v[92] = 10'b1100011111;
    16'b1001000010000001: out_v[92] = 10'b1101001101;
    16'b0001110011010000: out_v[92] = 10'b1011010001;
    16'b0000100010010000: out_v[92] = 10'b0011111110;
    16'b1001100011010001: out_v[92] = 10'b0011000101;
    16'b0001100010000000: out_v[92] = 10'b0100000001;
    16'b1001100000010000: out_v[92] = 10'b0001110111;
    16'b1001100010010001: out_v[92] = 10'b0111011111;
    16'b1001110010000000: out_v[92] = 10'b1111101111;
    16'b0000000010010001: out_v[92] = 10'b1111110001;
    16'b0000100000000001: out_v[92] = 10'b1011101001;
    16'b0001100010010000: out_v[92] = 10'b1010110011;
    16'b0000100010010001: out_v[92] = 10'b0111001100;
    16'b0000110010010001: out_v[92] = 10'b1100100110;
    16'b1001110011010001: out_v[92] = 10'b1000010101;
    16'b0001110010010001: out_v[92] = 10'b0101101100;
    16'b1000100010000001: out_v[92] = 10'b1000001001;
    16'b1001110000010000: out_v[92] = 10'b0100010101;
    16'b1001010000010000: out_v[92] = 10'b1000001011;
    16'b0000110010000000: out_v[92] = 10'b1100011001;
    16'b0001100010000001: out_v[92] = 10'b1111101010;
    16'b1001000010010000: out_v[92] = 10'b0011100000;
    16'b1001100010000000: out_v[92] = 10'b1101011001;
    16'b0001110010000001: out_v[92] = 10'b0110011111;
    16'b0000110010010000: out_v[92] = 10'b0000100110;
    16'b1001111011010000: out_v[92] = 10'b0010000111;
    16'b0001110011010001: out_v[92] = 10'b0010111111;
    16'b1001000010010001: out_v[92] = 10'b1001011111;
    16'b0001111001010011: out_v[92] = 10'b1010100110;
    16'b0000000001000000: out_v[92] = 10'b1001110111;
    16'b0000000001000010: out_v[92] = 10'b0010011111;
    16'b0000000000010010: out_v[92] = 10'b0101111001;
    16'b0000110001010011: out_v[92] = 10'b1111010111;
    16'b0000110000010011: out_v[92] = 10'b1111110000;
    16'b0001111000010011: out_v[92] = 10'b0001100100;
    16'b0000010001010010: out_v[92] = 10'b0111000010;
    16'b0000000001010010: out_v[92] = 10'b0011001111;
    16'b0000110001010010: out_v[92] = 10'b1111110110;
    16'b1001111000010011: out_v[92] = 10'b1000101101;
    16'b0000111001010011: out_v[92] = 10'b1111100011;
    16'b0000000000010011: out_v[92] = 10'b0100110001;
    16'b1001111001010011: out_v[92] = 10'b1010111111;
    16'b0000111000010011: out_v[92] = 10'b0110111100;
    16'b0001110000010011: out_v[92] = 10'b0110100001;
    16'b1001111000010010: out_v[92] = 10'b1110100010;
    16'b0000000000010000: out_v[92] = 10'b1111110100;
    16'b0000111001010010: out_v[92] = 10'b1101111010;
    16'b0000000001010011: out_v[92] = 10'b0101001100;
    16'b0000010001010011: out_v[92] = 10'b1111001101;
    16'b0000000000000010: out_v[92] = 10'b1011100110;
    16'b0000001001010010: out_v[92] = 10'b0010110010;
    16'b0000011001010010: out_v[92] = 10'b1010100111;
    16'b0001111000010010: out_v[92] = 10'b0111010111;
    16'b0000000000000000: out_v[92] = 10'b0111101001;
    16'b0000010000010011: out_v[92] = 10'b0111011011;
    16'b0000000001010000: out_v[92] = 10'b1000001111;
    16'b0001110001010011: out_v[92] = 10'b1011000000;
    16'b0000010000010010: out_v[92] = 10'b1000111100;
    16'b0000010001000010: out_v[92] = 10'b1100000111;
    16'b0000110000010010: out_v[92] = 10'b1110110100;
    16'b0000111000010000: out_v[92] = 10'b0010010101;
    16'b0000111000010010: out_v[92] = 10'b0000011100;
    16'b0001111000010001: out_v[92] = 10'b1100011110;
    16'b1001111000010001: out_v[92] = 10'b1110010000;
    16'b0000001000010000: out_v[92] = 10'b0111010010;
    16'b1001111000000001: out_v[92] = 10'b1010011101;
    16'b1101110010000001: out_v[92] = 10'b0110100110;
    16'b0000011000010000: out_v[92] = 10'b1010010101;
    16'b1001110000010010: out_v[92] = 10'b1100010100;
    16'b1001110000000001: out_v[92] = 10'b0010010101;
    16'b0001111000010000: out_v[92] = 10'b1011110100;
    16'b1001111000000011: out_v[92] = 10'b1111111010;
    16'b1000110010000011: out_v[92] = 10'b0100001010;
    16'b0000110001000010: out_v[92] = 10'b0010111111;
    16'b1001111010010011: out_v[92] = 10'b0000110101;
    16'b1001111010000011: out_v[92] = 10'b0011010011;
    16'b1001110010010010: out_v[92] = 10'b1110000110;
    16'b1001100010000011: out_v[92] = 10'b1010010110;
    16'b0000110001010000: out_v[92] = 10'b0110011101;
    16'b0000110000010000: out_v[92] = 10'b0011110110;
    16'b1001110010000011: out_v[92] = 10'b0011110110;
    16'b0000011000010010: out_v[92] = 10'b0001011101;
    16'b1101110010000011: out_v[92] = 10'b1110110101;
    16'b1001110000000011: out_v[92] = 10'b0110010110;
    16'b1000110010000001: out_v[92] = 10'b0000001011;
    16'b1001101000010010: out_v[92] = 10'b1011011011;
    16'b1001110010000010: out_v[92] = 10'b0100111000;
    16'b0000001001010000: out_v[92] = 10'b1001000000;
    16'b1001001000010010: out_v[92] = 10'b1000101011;
    16'b1001111001010000: out_v[92] = 10'b1101011010;
    16'b1000001001010000: out_v[92] = 10'b1101100001;
    16'b0000001000010010: out_v[92] = 10'b0101011001;
    16'b0000111001010000: out_v[92] = 10'b1000111001;
    16'b0001000001010010: out_v[92] = 10'b0110001111;
    16'b1001101000010011: out_v[92] = 10'b1111111111;
    16'b0000100001010000: out_v[92] = 10'b1001011001;
    16'b1000001001000000: out_v[92] = 10'b0010100011;
    16'b0000101001010000: out_v[92] = 10'b1111000000;
    16'b0001101001010000: out_v[92] = 10'b0111100011;
    16'b1000101001010000: out_v[92] = 10'b0101001110;
    16'b0001111001010001: out_v[92] = 10'b0110011100;
    16'b0000000001010001: out_v[92] = 10'b0111001001;
    16'b1001001000010011: out_v[92] = 10'b0011001010;
    16'b1001111001010010: out_v[92] = 10'b0100011010;
    16'b1001111001010001: out_v[92] = 10'b0010001001;
    16'b0001000001010001: out_v[92] = 10'b1110001100;
    16'b0001000001010000: out_v[92] = 10'b1000000101;
    16'b0000100001010010: out_v[92] = 10'b1010001011;
    16'b0000110001000000: out_v[92] = 10'b1100011011;
    16'b0000100001000000: out_v[92] = 10'b0110001011;
    16'b0001001001010001: out_v[92] = 10'b1100000111;
    16'b0001001000010010: out_v[92] = 10'b0101001100;
    16'b0001001000010011: out_v[92] = 10'b0111011011;
    16'b1001001001010000: out_v[92] = 10'b0011100011;
    16'b1001101001010001: out_v[92] = 10'b0111001111;
    16'b1001001010000011: out_v[92] = 10'b1000101011;
    16'b1001101001010000: out_v[92] = 10'b1111100110;
    16'b1001001001010001: out_v[92] = 10'b0101111110;
    16'b1000111001010000: out_v[92] = 10'b0111001010;
    16'b1000101001000000: out_v[92] = 10'b0000110101;
    16'b0001001000010000: out_v[92] = 10'b0011010110;
    16'b0001101001010001: out_v[92] = 10'b0001001010;
    16'b0001001001010010: out_v[92] = 10'b0011011000;
    16'b1001000010000000: out_v[92] = 10'b0000110111;
    16'b1001000010000010: out_v[92] = 10'b1001010001;
    16'b1001001000010000: out_v[92] = 10'b0111110110;
    16'b1001001000000010: out_v[92] = 10'b0000111101;
    16'b0000001000010001: out_v[92] = 10'b0111110011;
    16'b1001111000000010: out_v[92] = 10'b0111010001;
    16'b1001001010000010: out_v[92] = 10'b0001111111;
    16'b1001001000000011: out_v[92] = 10'b1011001111;
    16'b1001001000010001: out_v[92] = 10'b0101010101;
    16'b0000001000010011: out_v[92] = 10'b1101001001;
    16'b1000001000010010: out_v[92] = 10'b0111010001;
    16'b1001000000000010: out_v[92] = 10'b1100011011;
    16'b1000000010000010: out_v[92] = 10'b1100010001;
    16'b1001001010010010: out_v[92] = 10'b1100011011;
    16'b1001000000000000: out_v[92] = 10'b0110011000;
    16'b1001000000000011: out_v[92] = 10'b0111000110;
    16'b1001000000000001: out_v[92] = 10'b0101010111;
    16'b1001001000000000: out_v[92] = 10'b0000010011;
    16'b1000000010000000: out_v[92] = 10'b1010010010;
    16'b1001010010000000: out_v[92] = 10'b0010110010;
    16'b1001000000010010: out_v[92] = 10'b1101011111;
    16'b1001011000010000: out_v[92] = 10'b1000011110;
    16'b0001001000010001: out_v[92] = 10'b0000011011;
    16'b1001111010000010: out_v[92] = 10'b1011110110;
    16'b1001001010000000: out_v[92] = 10'b1001010011;
    16'b0000101001000001: out_v[92] = 10'b1011110111;
    16'b0001110000010010: out_v[92] = 10'b0010010010;
    16'b0000000000000011: out_v[92] = 10'b0010100111;
    16'b0000100000010000: out_v[92] = 10'b1011001010;
    16'b0000100000000011: out_v[92] = 10'b0011100010;
    16'b0000110000000000: out_v[92] = 10'b0010111010;
    16'b0000100000010010: out_v[92] = 10'b0010111010;
    16'b1000111001000000: out_v[92] = 10'b0011110010;
    16'b1000101001000001: out_v[92] = 10'b1010110010;
    16'b0001000000010000: out_v[92] = 10'b0000100000;
    16'b1000111001000001: out_v[92] = 10'b1011100110;
    16'b0001110001010000: out_v[92] = 10'b0110110000;
    16'b0000111001000001: out_v[92] = 10'b0010110010;
    16'b0000110000000001: out_v[92] = 10'b1001111110;
    16'b0001100001010000: out_v[92] = 10'b1110101111;
    16'b0000110000000011: out_v[92] = 10'b1011011001;
    16'b0000110001000001: out_v[92] = 10'b1010110100;
    16'b0001100001010010: out_v[92] = 10'b0011001101;
    16'b1000001001000001: out_v[92] = 10'b0111110100;
    16'b0001000000010010: out_v[92] = 10'b1101100000;
    16'b0000100000000000: out_v[92] = 10'b0010111010;
    16'b0001100000010010: out_v[92] = 10'b0001100001;
    16'b0001110000010000: out_v[92] = 10'b0001101000;
    16'b1000101000000001: out_v[92] = 10'b0011100100;
    16'b0001110001010010: out_v[92] = 10'b1111010100;
    16'b0000100000010011: out_v[92] = 10'b1010110110;
    16'b0000100001000001: out_v[92] = 10'b1011100100;
    16'b0000100000000010: out_v[92] = 10'b1010101110;
    16'b1000001000000001: out_v[92] = 10'b0010110110;
    16'b0001100000010000: out_v[92] = 10'b0101011011;
    16'b1000110000000010: out_v[92] = 10'b1101111011;
    16'b1000111010000010: out_v[92] = 10'b0110111010;
    16'b1001011010000010: out_v[92] = 10'b0111100011;
    16'b1000111000000010: out_v[92] = 10'b1011100001;
    16'b1000010000000000: out_v[92] = 10'b1101101010;
    16'b1000111000000000: out_v[92] = 10'b0111100010;
    16'b0000010000000000: out_v[92] = 10'b0001001010;
    16'b1000011000000010: out_v[92] = 10'b1011101011;
    16'b1000110000000011: out_v[92] = 10'b1111011001;
    16'b0000110000000010: out_v[92] = 10'b1001001010;
    16'b0000110001000011: out_v[92] = 10'b0110010001;
    16'b1000011000000000: out_v[92] = 10'b0011101010;
    16'b1000110000000000: out_v[92] = 10'b1010101010;
    16'b1000111010000000: out_v[92] = 10'b1011110000;
    16'b0000010000000001: out_v[92] = 10'b1011000011;
    16'b0000110000001001: out_v[92] = 10'b1100011011;
    16'b1001011010000000: out_v[92] = 10'b1011000110;
    16'b0000010000000010: out_v[92] = 10'b1000101110;
    16'b1001111010000000: out_v[92] = 10'b1011011010;
    16'b0000110001010001: out_v[92] = 10'b1101001100;
    16'b0000010000000011: out_v[92] = 10'b0001100101;
    16'b1000110010000000: out_v[92] = 10'b1111001010;
    16'b1000010000000010: out_v[92] = 10'b1110010001;
    16'b0000110000001000: out_v[92] = 10'b0010111010;
    16'b1000111000000011: out_v[92] = 10'b1011011111;
    16'b1001000011010000: out_v[92] = 10'b0111100011;
    16'b1001001010010000: out_v[92] = 10'b1010000101;
    16'b1001000000010000: out_v[92] = 10'b1011000100;
    16'b1001001011010000: out_v[92] = 10'b0110000000;
    16'b1001001011000000: out_v[92] = 10'b0110000111;
    16'b1001000001010000: out_v[92] = 10'b1101000111;
    16'b1001111010010010: out_v[92] = 10'b0111011101;
    16'b1000001000010000: out_v[92] = 10'b1101111011;
    16'b0001000010010000: out_v[92] = 10'b1011100110;
    16'b1001111011010010: out_v[92] = 10'b1111001001;
    16'b0001111001010010: out_v[92] = 10'b1101010101;
    16'b1001111001000011: out_v[92] = 10'b1110000001;
    16'b0001011000010010: out_v[92] = 10'b1110110101;
    16'b1001011000000010: out_v[92] = 10'b0011001111;
    16'b1001111011000011: out_v[92] = 10'b1011001010;
    16'b1001111011000010: out_v[92] = 10'b0111001000;
    16'b1001111011010011: out_v[92] = 10'b1111011001;
    16'b0001111000000011: out_v[92] = 10'b1101010111;
    16'b1001011000010010: out_v[92] = 10'b0101011110;
    16'b1001001001010010: out_v[92] = 10'b0010011100;
    16'b0000001000000010: out_v[92] = 10'b1100001101;
    16'b1001000010010010: out_v[92] = 10'b1000101010;
    16'b1001001011010010: out_v[92] = 10'b1000100110;
    16'b0000001000000000: out_v[92] = 10'b1100110101;
    16'b1001010010010000: out_v[92] = 10'b1000011111;
    default: out_v[92] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000010000000000: out_v[93] = 10'b1001100000;
    16'b1000010010000000: out_v[93] = 10'b0111011100;
    16'b0000100000000000: out_v[93] = 10'b0011000111;
    16'b0000110000000000: out_v[93] = 10'b1101010001;
    16'b1000110000000000: out_v[93] = 10'b0011001011;
    16'b0000000000000000: out_v[93] = 10'b1010100010;
    16'b0000110010000001: out_v[93] = 10'b0011100101;
    16'b1000010000000000: out_v[93] = 10'b0000010111;
    16'b0010110000000000: out_v[93] = 10'b0001011010;
    16'b0000100010000000: out_v[93] = 10'b0100111001;
    16'b0000110010100000: out_v[93] = 10'b1111011011;
    16'b0000010010000001: out_v[93] = 10'b0101011000;
    16'b0000010010000000: out_v[93] = 10'b1010101010;
    16'b0000110010100001: out_v[93] = 10'b0110011001;
    16'b0000010010100000: out_v[93] = 10'b1100101000;
    16'b0010010000000000: out_v[93] = 10'b0000010000;
    16'b0000010010100001: out_v[93] = 10'b1100100010;
    16'b0000110010000000: out_v[93] = 10'b0011000101;
    16'b0000100010000001: out_v[93] = 10'b0110110100;
    16'b0010010010000000: out_v[93] = 10'b0011110101;
    16'b0000000010000000: out_v[93] = 10'b0010001001;
    16'b0000000010000001: out_v[93] = 10'b0011010101;
    16'b1000110010000000: out_v[93] = 10'b0000101111;
    16'b0000000000100000: out_v[93] = 10'b0110010010;
    16'b0000000010100001: out_v[93] = 10'b0101001100;
    16'b0000101010000001: out_v[93] = 10'b1001111100;
    16'b0000100001000000: out_v[93] = 10'b0011011110;
    16'b0000100010100001: out_v[93] = 10'b1110110110;
    16'b0000000011000001: out_v[93] = 10'b1110110011;
    16'b0000100000000001: out_v[93] = 10'b0111100110;
    16'b1000100010000000: out_v[93] = 10'b1011011010;
    16'b1000100011000001: out_v[93] = 10'b1110101011;
    16'b1000100010000001: out_v[93] = 10'b0111001001;
    16'b0000100011000000: out_v[93] = 10'b1001011110;
    16'b0000100011000001: out_v[93] = 10'b0110110110;
    16'b1000100000000000: out_v[93] = 10'b0000100000;
    16'b0000101010100001: out_v[93] = 10'b1011110111;
    16'b0000000001000000: out_v[93] = 10'b1101001111;
    16'b0000100010100000: out_v[93] = 10'b0001111110;
    16'b0000000000000001: out_v[93] = 10'b0001001100;
    16'b1000000000000000: out_v[93] = 10'b1001101101;
    16'b0000001010000001: out_v[93] = 10'b0010010101;
    16'b0000100000100000: out_v[93] = 10'b1001001000;
    16'b0000000010100000: out_v[93] = 10'b1111001001;
    16'b0000100001000001: out_v[93] = 10'b1010101011;
    16'b1000000010000000: out_v[93] = 10'b0001110111;
    16'b1000000010000001: out_v[93] = 10'b0000100110;
    16'b0000010000100000: out_v[93] = 10'b0010110000;
    16'b0010100000000000: out_v[93] = 10'b0110100001;
    16'b0010000000000000: out_v[93] = 10'b0100110101;
    16'b0010000010000000: out_v[93] = 10'b1111000010;
    16'b0000000011000000: out_v[93] = 10'b0001111010;
    16'b0000110011000000: out_v[93] = 10'b0001001001;
    16'b0000110011000001: out_v[93] = 10'b0001101011;
    16'b0000110001000000: out_v[93] = 10'b0011100000;
    16'b0010100010000001: out_v[93] = 10'b1111000010;
    16'b0010100010000000: out_v[93] = 10'b1100101011;
    default: out_v[93] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000001010000000: out_v[94] = 10'b0110001011;
    16'b0100001010000000: out_v[94] = 10'b1000101011;
    16'b0100001110101000: out_v[94] = 10'b1101100111;
    16'b0000000010000000: out_v[94] = 10'b1001101010;
    16'b0000001000000000: out_v[94] = 10'b1110110010;
    16'b0000001110101010: out_v[94] = 10'b0100010001;
    16'b0100000110101000: out_v[94] = 10'b0010011011;
    16'b0000001100101000: out_v[94] = 10'b1010111011;
    16'b0000000110101000: out_v[94] = 10'b0110001010;
    16'b0100000010000000: out_v[94] = 10'b1000101100;
    16'b0100001010101000: out_v[94] = 10'b1011110111;
    16'b0100000010101000: out_v[94] = 10'b0101011110;
    16'b0100000010100000: out_v[94] = 10'b1101111110;
    16'b0000001010100000: out_v[94] = 10'b1100000001;
    16'b0100001000001000: out_v[94] = 10'b1100010111;
    16'b0100001010100000: out_v[94] = 10'b0000011011;
    16'b0100000000000000: out_v[94] = 10'b1100101111;
    16'b0000001110101000: out_v[94] = 10'b1110010001;
    16'b0000001010101000: out_v[94] = 10'b1100101100;
    16'b0100001000000000: out_v[94] = 10'b0011100001;
    16'b0000000010101000: out_v[94] = 10'b1110110111;
    16'b0100001000000001: out_v[94] = 10'b1000011100;
    16'b0100000110101010: out_v[94] = 10'b1111100100;
    16'b0000000010100000: out_v[94] = 10'b0100110001;
    16'b0100000000000001: out_v[94] = 10'b0110101001;
    16'b0000000100101000: out_v[94] = 10'b0111000001;
    16'b0100001110001000: out_v[94] = 10'b0000011011;
    16'b0100001010001000: out_v[94] = 10'b1111001110;
    16'b0000000000000000: out_v[94] = 10'b1111011000;
    16'b0100001110101010: out_v[94] = 10'b0110011011;
    16'b0100001110101001: out_v[94] = 10'b0001011001;
    16'b0100000110001000: out_v[94] = 10'b0011001111;
    16'b0100000010001000: out_v[94] = 10'b0110010110;
    16'b0100001100101000: out_v[94] = 10'b1100100110;
    16'b0100001010000001: out_v[94] = 10'b0000001100;
    16'b0000000110101010: out_v[94] = 10'b1011100110;
    16'b0000001010000010: out_v[94] = 10'b1011110101;
    16'b1000001010000000: out_v[94] = 10'b0111110111;
    16'b0000001000000010: out_v[94] = 10'b0101100110;
    16'b1000001000000000: out_v[94] = 10'b1100110110;
    16'b0100001000100000: out_v[94] = 10'b1001010111;
    16'b1000001000000010: out_v[94] = 10'b0111101110;
    16'b1100001000000000: out_v[94] = 10'b0111000100;
    16'b0100001100000010: out_v[94] = 10'b1001101011;
    16'b0000001000100000: out_v[94] = 10'b1110100000;
    16'b1000000000000010: out_v[94] = 10'b1110010101;
    16'b0100001100000000: out_v[94] = 10'b1011001101;
    16'b0000000100100010: out_v[94] = 10'b1101100101;
    16'b1100001000000010: out_v[94] = 10'b1111011011;
    16'b0000000100000010: out_v[94] = 10'b0101101101;
    16'b0000001100000010: out_v[94] = 10'b1011100011;
    16'b0100000010000001: out_v[94] = 10'b1111100100;
    16'b0000000100000000: out_v[94] = 10'b0000000111;
    16'b0000000000000010: out_v[94] = 10'b1010000100;
    16'b1000001010000010: out_v[94] = 10'b1110110111;
    16'b0000001100000000: out_v[94] = 10'b1100110000;
    16'b1000001000100010: out_v[94] = 10'b0010101100;
    16'b0100001000000010: out_v[94] = 10'b1110111101;
    16'b0001000010000000: out_v[94] = 10'b0111100000;
    16'b0000000110000000: out_v[94] = 10'b1101011001;
    16'b0000001010000001: out_v[94] = 10'b1101001011;
    16'b0001001010000000: out_v[94] = 10'b0001010110;
    16'b0100001010100001: out_v[94] = 10'b1010100010;
    16'b0000000000100000: out_v[94] = 10'b0010111000;
    16'b0000001100100000: out_v[94] = 10'b0011011110;
    16'b0000001000101000: out_v[94] = 10'b1011011011;
    16'b0000001100001000: out_v[94] = 10'b1101011111;
    16'b0000000000001000: out_v[94] = 10'b1010100111;
    16'b0000001000001000: out_v[94] = 10'b0100110111;
    16'b0100000010100001: out_v[94] = 10'b0111101010;
    16'b0000000110100000: out_v[94] = 10'b0011100000;
    16'b0000010010000000: out_v[94] = 10'b0010101101;
    16'b0000000101101000: out_v[94] = 10'b1111001111;
    16'b0000000100101010: out_v[94] = 10'b0111101001;
    16'b0000000100100000: out_v[94] = 10'b0001010110;
    16'b0000010000000000: out_v[94] = 10'b0111101011;
    16'b0000000110001000: out_v[94] = 10'b1011011001;
    16'b0000000100001000: out_v[94] = 10'b0111000111;
    16'b0000000000101000: out_v[94] = 10'b0101101110;
    default: out_v[94] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010000000000010: out_v[95] = 10'b0101101101;
    16'b0011000001000010: out_v[95] = 10'b1101100011;
    16'b0010000000000000: out_v[95] = 10'b0001000111;
    16'b0000000000000000: out_v[95] = 10'b0011001111;
    16'b0010000001000000: out_v[95] = 10'b0000010000;
    16'b0000000001000000: out_v[95] = 10'b0001000111;
    16'b0011000000000000: out_v[95] = 10'b1111000010;
    16'b0001000000000000: out_v[95] = 10'b0101001011;
    16'b0000000000000010: out_v[95] = 10'b0110010110;
    16'b0010000000001010: out_v[95] = 10'b1110011010;
    16'b0010000000001000: out_v[95] = 10'b0001010001;
    16'b0010000000000001: out_v[95] = 10'b1001001111;
    16'b0000000000000001: out_v[95] = 10'b1000110100;
    16'b0010000001000010: out_v[95] = 10'b0000010111;
    16'b0001000000000001: out_v[95] = 10'b0100110011;
    16'b0000000000001000: out_v[95] = 10'b1100000111;
    16'b0011000000000010: out_v[95] = 10'b0101101000;
    16'b0011000001000000: out_v[95] = 10'b1111011011;
    16'b0011000000000001: out_v[95] = 10'b0011000100;
    16'b0011000000001000: out_v[95] = 10'b1010101011;
    16'b0010000001000001: out_v[95] = 10'b0110111111;
    16'b0001000000000010: out_v[95] = 10'b1101010000;
    16'b0011000010000000: out_v[95] = 10'b0011101010;
    16'b0000000010000000: out_v[95] = 10'b1000111110;
    16'b0001000001000000: out_v[95] = 10'b0000110101;
    16'b0011001010000000: out_v[95] = 10'b0101000110;
    16'b0010000000000100: out_v[95] = 10'b0110011100;
    16'b0000001010000000: out_v[95] = 10'b1100101110;
    16'b0111000010000100: out_v[95] = 10'b0111000110;
    16'b0010000010000000: out_v[95] = 10'b0100000110;
    16'b0001001010000000: out_v[95] = 10'b1011100011;
    16'b0001001000000000: out_v[95] = 10'b1111100011;
    16'b0010001010000000: out_v[95] = 10'b0000001110;
    16'b0110000000000100: out_v[95] = 10'b1110010111;
    16'b0111000000000100: out_v[95] = 10'b1110011100;
    16'b0000001000000000: out_v[95] = 10'b0001000101;
    16'b0000000000000100: out_v[95] = 10'b0111001001;
    16'b0001000010000000: out_v[95] = 10'b1100010101;
    16'b0100000000000100: out_v[95] = 10'b0010011010;
    16'b0011100000000010: out_v[95] = 10'b0001011110;
    16'b0111000000000110: out_v[95] = 10'b1001001001;
    16'b0011000000000110: out_v[95] = 10'b0100011000;
    16'b0101000000000110: out_v[95] = 10'b1101100010;
    16'b0011000000000100: out_v[95] = 10'b1110100010;
    16'b0001000000000011: out_v[95] = 10'b0010001100;
    16'b0000000000000011: out_v[95] = 10'b1101010110;
    16'b0011000000000011: out_v[95] = 10'b1100100011;
    16'b0010000000000011: out_v[95] = 10'b1010001100;
    16'b0000100000000100: out_v[95] = 10'b0011010011;
    16'b0000010000000010: out_v[95] = 10'b0111010111;
    16'b0110000000000110: out_v[95] = 10'b0111010101;
    16'b0000010000000000: out_v[95] = 10'b1000101110;
    16'b0000100000000000: out_v[95] = 10'b1011110000;
    16'b0010000000000110: out_v[95] = 10'b1101110110;
    16'b0000000000000110: out_v[95] = 10'b0011101010;
    16'b0100000000000110: out_v[95] = 10'b1110001011;
    16'b0001010000000010: out_v[95] = 10'b1100100011;
    16'b0000010000000110: out_v[95] = 10'b1100111110;
    16'b0001100000000000: out_v[95] = 10'b1000100000;
    16'b0100010000000110: out_v[95] = 10'b1101001100;
    default: out_v[95] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000110000100000: out_v[96] = 10'b0101010110;
    16'b0000000000100010: out_v[96] = 10'b1000100101;
    16'b0000100101100110: out_v[96] = 10'b0111011110;
    16'b0000100001100110: out_v[96] = 10'b0010111110;
    16'b0000100000100000: out_v[96] = 10'b1111010011;
    16'b0000100101000100: out_v[96] = 10'b0111011011;
    16'b0000000000000110: out_v[96] = 10'b1011010101;
    16'b0000100001000100: out_v[96] = 10'b1100110101;
    16'b0000010000100110: out_v[96] = 10'b1111110011;
    16'b0000010000000000: out_v[96] = 10'b0010011101;
    16'b0000100000110010: out_v[96] = 10'b1101001011;
    16'b0000000001100110: out_v[96] = 10'b1111110111;
    16'b1000100000110000: out_v[96] = 10'b1001011101;
    16'b0000100000110110: out_v[96] = 10'b0110011011;
    16'b0000100000000000: out_v[96] = 10'b0011110110;
    16'b0000110000000100: out_v[96] = 10'b0010101111;
    16'b0000110000100100: out_v[96] = 10'b1000010011;
    16'b0000110000000000: out_v[96] = 10'b0111001011;
    16'b0000100001100100: out_v[96] = 10'b0111110011;
    16'b0000110001100110: out_v[96] = 10'b1111111101;
    16'b0000100000000010: out_v[96] = 10'b0010011011;
    16'b0000100000100010: out_v[96] = 10'b0111000101;
    16'b0000110101100100: out_v[96] = 10'b0001010111;
    16'b0000110000100110: out_v[96] = 10'b1111011100;
    16'b0000100000000100: out_v[96] = 10'b1011110110;
    16'b0000110101000100: out_v[96] = 10'b0111010010;
    16'b0000000000010000: out_v[96] = 10'b1001011100;
    16'b0100100000100010: out_v[96] = 10'b1011001101;
    16'b0000100101100100: out_v[96] = 10'b1111101111;
    16'b0000100000100110: out_v[96] = 10'b0011011110;
    16'b0000000000100000: out_v[96] = 10'b0100011101;
    16'b0000010101100110: out_v[96] = 10'b1101110111;
    16'b0000100000110000: out_v[96] = 10'b1011010100;
    16'b0000110001100100: out_v[96] = 10'b0011011111;
    16'b0000110100000100: out_v[96] = 10'b1010011001;
    16'b0000000001100010: out_v[96] = 10'b1011001010;
    16'b0000110101100110: out_v[96] = 10'b0110010011;
    16'b0000100001100010: out_v[96] = 10'b1011011000;
    16'b0000000101100110: out_v[96] = 10'b0101111110;
    16'b0000010000000100: out_v[96] = 10'b0010110011;
    16'b0000000000000000: out_v[96] = 10'b0011000011;
    16'b0000100000100100: out_v[96] = 10'b1111011100;
    16'b1000100000110010: out_v[96] = 10'b1001001111;
    16'b0100100000110010: out_v[96] = 10'b0011011110;
    16'b0000000000100110: out_v[96] = 10'b1100110110;
    16'b0000010001100110: out_v[96] = 10'b1110010011;
    16'b0000110100100100: out_v[96] = 10'b0101001011;
    16'b0000000000110010: out_v[96] = 10'b0000100010;
    16'b1100000000110000: out_v[96] = 10'b0100000001;
    16'b1000000000110000: out_v[96] = 10'b0001011011;
    16'b1000000000010000: out_v[96] = 10'b0000111111;
    16'b1000010000010000: out_v[96] = 10'b0010010011;
    16'b1000000000000000: out_v[96] = 10'b0111100110;
    16'b0000000000110000: out_v[96] = 10'b1100011111;
    16'b0100000000110000: out_v[96] = 10'b0010101111;
    16'b1100000000110010: out_v[96] = 10'b1110010000;
    16'b1000000000100000: out_v[96] = 10'b0111110000;
    16'b0100000000110010: out_v[96] = 10'b1001001110;
    16'b1000000000110010: out_v[96] = 10'b1101100001;
    16'b1100100000110010: out_v[96] = 10'b0100110011;
    16'b0000000000010100: out_v[96] = 10'b0100001100;
    16'b1000000000110100: out_v[96] = 10'b0010110011;
    16'b1000001000000100: out_v[96] = 10'b1011011010;
    16'b1000001000100000: out_v[96] = 10'b1001011000;
    16'b1000010000000000: out_v[96] = 10'b1100011100;
    16'b1000000000000100: out_v[96] = 10'b0111000110;
    16'b1000000100010100: out_v[96] = 10'b1001100110;
    16'b1000001000000000: out_v[96] = 10'b0100000010;
    16'b1000001000100100: out_v[96] = 10'b0110011011;
    16'b0000010000010000: out_v[96] = 10'b1100001000;
    16'b1000100000100000: out_v[96] = 10'b1000100110;
    16'b1000000000100100: out_v[96] = 10'b1011011010;
    16'b1000100000100100: out_v[96] = 10'b1101010111;
    16'b1000000000010100: out_v[96] = 10'b1010100110;
    16'b1000000100000000: out_v[96] = 10'b0001111101;
    16'b1000000100000100: out_v[96] = 10'b1001000100;
    16'b1000101000100100: out_v[96] = 10'b1110111111;
    16'b1100101000000010: out_v[96] = 10'b1110010100;
    16'b1000100000100010: out_v[96] = 10'b0111001100;
    16'b1000010000100000: out_v[96] = 10'b1101000110;
    16'b1000100000100110: out_v[96] = 10'b0111110110;
    16'b1000110000100010: out_v[96] = 10'b0101001111;
    16'b1000100000110100: out_v[96] = 10'b1010011100;
    16'b1100100000000010: out_v[96] = 10'b1011011101;
    16'b1000101000100000: out_v[96] = 10'b1110011100;
    16'b1000110000100000: out_v[96] = 10'b1010001110;
    16'b1000001000010100: out_v[96] = 10'b1000110101;
    16'b1000101000100010: out_v[96] = 10'b1110110011;
    16'b1000100000000000: out_v[96] = 10'b0011100010;
    16'b1000100000000100: out_v[96] = 10'b0001010110;
    16'b1100100000100010: out_v[96] = 10'b1001011010;
    16'b0000010100010000: out_v[96] = 10'b1100010100;
    16'b0000001000110000: out_v[96] = 10'b1110001100;
    16'b0000010000010100: out_v[96] = 10'b0100001000;
    16'b0000000000110100: out_v[96] = 10'b0101011100;
    16'b1000010000010100: out_v[96] = 10'b0101010000;
    16'b0000100000110100: out_v[96] = 10'b0110011001;
    16'b0000010100010100: out_v[96] = 10'b0110111010;
    16'b0000010000110000: out_v[96] = 10'b0011010110;
    16'b0000010000110100: out_v[96] = 10'b1011011110;
    16'b0000110000110010: out_v[96] = 10'b0101111011;
    16'b0000100000010010: out_v[96] = 10'b1010011010;
    16'b0000110000110110: out_v[96] = 10'b1011011010;
    16'b0000000100010100: out_v[96] = 10'b0100001010;
    16'b0000000000000100: out_v[96] = 10'b1000001011;
    16'b0000110000110100: out_v[96] = 10'b0000001011;
    16'b0000110000110000: out_v[96] = 10'b0110011101;
    16'b1000010000110000: out_v[96] = 10'b1110001100;
    16'b1000100000010010: out_v[96] = 10'b0000011011;
    16'b1000100000010000: out_v[96] = 10'b1100110000;
    16'b1000000000100010: out_v[96] = 10'b1100100110;
    16'b1000100000000010: out_v[96] = 10'b0011010010;
    16'b1000110000000010: out_v[96] = 10'b0110011000;
    16'b1000110000000000: out_v[96] = 10'b0001111100;
    16'b1000100001000010: out_v[96] = 10'b0100111100;
    16'b1000100001000000: out_v[96] = 10'b0000011011;
    16'b1100000000100000: out_v[96] = 10'b1000111010;
    16'b1000100001010010: out_v[96] = 10'b1111010011;
    16'b0000010000100000: out_v[96] = 10'b0011111011;
    16'b0000010000110110: out_v[96] = 10'b1001100111;
    16'b0000100000010000: out_v[96] = 10'b1111100010;
    16'b1000010000110010: out_v[96] = 10'b1110100000;
    16'b1000000000010010: out_v[96] = 10'b1101000001;
    16'b0100000000010000: out_v[96] = 10'b0011010010;
    16'b0000010000100010: out_v[96] = 10'b1000110110;
    16'b0000010000110010: out_v[96] = 10'b1010110010;
    16'b1000000000000010: out_v[96] = 10'b0101000111;
    16'b0000000000010010: out_v[96] = 10'b0101110010;
    16'b1000010000100010: out_v[96] = 10'b1110000010;
    16'b0000000000110110: out_v[96] = 10'b1110100001;
    16'b0100010000010000: out_v[96] = 10'b1010111111;
    16'b0000010100110110: out_v[96] = 10'b0111110100;
    16'b0100010000010100: out_v[96] = 10'b1000001111;
    16'b0000001000000100: out_v[96] = 10'b0011110010;
    16'b0000001000000000: out_v[96] = 10'b0001000011;
    16'b1010001000000100: out_v[96] = 10'b1100001011;
    16'b1000100100010100: out_v[96] = 10'b1111101010;
    16'b1010001000010000: out_v[96] = 10'b0011000011;
    16'b1100000000000000: out_v[96] = 10'b1001011100;
    16'b1000001000010000: out_v[96] = 10'b1011100101;
    16'b0010001000000100: out_v[96] = 10'b1011000111;
    16'b1100000000010000: out_v[96] = 10'b1011111000;
    16'b1010001000000000: out_v[96] = 10'b1010101101;
    16'b1010001000010100: out_v[96] = 10'b1100000111;
    16'b0000001000010000: out_v[96] = 10'b1011101100;
    16'b1000100000010100: out_v[96] = 10'b1011110011;
    16'b0010001000010100: out_v[96] = 10'b1111101000;
    16'b0010001000000000: out_v[96] = 10'b1011110010;
    16'b0000001000010100: out_v[96] = 10'b1111000110;
    16'b0000100000010100: out_v[96] = 10'b0001011000;
    16'b0010001000010000: out_v[96] = 10'b0010110001;
    16'b1000100100100010: out_v[96] = 10'b0111010001;
    16'b1000100100100000: out_v[96] = 10'b0010100110;
    16'b0000010100000000: out_v[96] = 10'b0111110101;
    16'b1000000100100000: out_v[96] = 10'b1010100100;
    16'b0000000100000000: out_v[96] = 10'b1011100001;
    16'b1000100100000000: out_v[96] = 10'b0010101111;
    16'b1000010100000000: out_v[96] = 10'b0100101110;
    16'b0000110100000000: out_v[96] = 10'b0110101110;
    16'b0000100100000000: out_v[96] = 10'b0110000101;
    16'b0001110110000000: out_v[96] = 10'b1101101101;
    16'b1000100100000010: out_v[96] = 10'b0011111011;
    16'b1000110000110000: out_v[96] = 10'b0110011000;
    16'b1000110000010000: out_v[96] = 10'b1101100010;
    16'b1000110000110010: out_v[96] = 10'b1000000101;
    16'b0000110000010000: out_v[96] = 10'b1111110110;
    16'b1100100000010010: out_v[96] = 10'b0110100101;
    16'b1000110000010010: out_v[96] = 10'b1110001111;
    default: out_v[96] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000010000000000: out_v[97] = 10'b0100111111;
    16'b0001010000001000: out_v[97] = 10'b1111100000;
    16'b0101010000011101: out_v[97] = 10'b0100111111;
    16'b0000000010000000: out_v[97] = 10'b1011010101;
    16'b0000010000000101: out_v[97] = 10'b1000011000;
    16'b1101010000011101: out_v[97] = 10'b1001100001;
    16'b1000000000000100: out_v[97] = 10'b1111010011;
    16'b0101010000001001: out_v[97] = 10'b1010101011;
    16'b1000000000010101: out_v[97] = 10'b1101100111;
    16'b0000010010000000: out_v[97] = 10'b0101011010;
    16'b0101010000011001: out_v[97] = 10'b0101011111;
    16'b0000010000001000: out_v[97] = 10'b1101000001;
    16'b0101000010010001: out_v[97] = 10'b1011010101;
    16'b0000010000010101: out_v[97] = 10'b1100001001;
    16'b0101010000010001: out_v[97] = 10'b1111001010;
    16'b0101000010001001: out_v[97] = 10'b0110110001;
    16'b1000010000010101: out_v[97] = 10'b0011001011;
    16'b0000010000010001: out_v[97] = 10'b1111011011;
    16'b1001010000010101: out_v[97] = 10'b1111110110;
    16'b0000000000000000: out_v[97] = 10'b0111111001;
    16'b0000000000000100: out_v[97] = 10'b1100100111;
    16'b0001010000001001: out_v[97] = 10'b0010011111;
    16'b0001000010001000: out_v[97] = 10'b0110010011;
    16'b0101000000001001: out_v[97] = 10'b1111011000;
    16'b0000000010001000: out_v[97] = 10'b1110011000;
    16'b0000000000001000: out_v[97] = 10'b0000111110;
    16'b0101000000011001: out_v[97] = 10'b1101001011;
    16'b0000010010010101: out_v[97] = 10'b0111011011;
    16'b0101000010011001: out_v[97] = 10'b0000010111;
    16'b0000000010010001: out_v[97] = 10'b0001111100;
    16'b1000010010010101: out_v[97] = 10'b1111111010;
    16'b0001010000011001: out_v[97] = 10'b1001111100;
    16'b0000000000010101: out_v[97] = 10'b0100100111;
    16'b0101000000011101: out_v[97] = 10'b0101010101;
    16'b0000010010000100: out_v[97] = 10'b0011000001;
    16'b0101000010000001: out_v[97] = 10'b1011010110;
    16'b0101010010011001: out_v[97] = 10'b0111011100;
    16'b0001000000001000: out_v[97] = 10'b1111100111;
    16'b0000010010001000: out_v[97] = 10'b0000011101;
    16'b0000010000000001: out_v[97] = 10'b1010111000;
    16'b0001010000010101: out_v[97] = 10'b0001111110;
    16'b0000010000000100: out_v[97] = 10'b0111001010;
    16'b0101010010011101: out_v[97] = 10'b1111110011;
    16'b1000010000000100: out_v[97] = 10'b1101001010;
    16'b0101010000010101: out_v[97] = 10'b1011111010;
    16'b0101010010010101: out_v[97] = 10'b1011110011;
    16'b0000000000000101: out_v[97] = 10'b0001101110;
    16'b0101000000000000: out_v[97] = 10'b0101011011;
    16'b0000000010000001: out_v[97] = 10'b0011011010;
    16'b0001000010000000: out_v[97] = 10'b0101011010;
    16'b0101000010010101: out_v[97] = 10'b1001000110;
    16'b0001010010001000: out_v[97] = 10'b1001001110;
    16'b0101010010001000: out_v[97] = 10'b1110001010;
    16'b0000010010010001: out_v[97] = 10'b1000110110;
    16'b0101010010010001: out_v[97] = 10'b0010111101;
    16'b0001010010000000: out_v[97] = 10'b0011010011;
    16'b0001000010000100: out_v[97] = 10'b1001101110;
    16'b0000000010000100: out_v[97] = 10'b1100110110;
    16'b0101010010000001: out_v[97] = 10'b0011100100;
    16'b0101000010000101: out_v[97] = 10'b1011111111;
    16'b0000010010000001: out_v[97] = 10'b1010111011;
    16'b0101000010001000: out_v[97] = 10'b0110111000;
    16'b0101000010000000: out_v[97] = 10'b1100011111;
    16'b0001000010010001: out_v[97] = 10'b1111001011;
    16'b0101010010000000: out_v[97] = 10'b0111110010;
    16'b0101010010001001: out_v[97] = 10'b1101010101;
    16'b0000000010010101: out_v[97] = 10'b1110111011;
    16'b0101010000001000: out_v[97] = 10'b0111011100;
    16'b0101010000000000: out_v[97] = 10'b0000110100;
    16'b0100010000001000: out_v[97] = 10'b0110010111;
    16'b0101010000000001: out_v[97] = 10'b1000001011;
    16'b0101000000001000: out_v[97] = 10'b1011101010;
    16'b0001010000000000: out_v[97] = 10'b0100011011;
    16'b0000000000010001: out_v[97] = 10'b1110110000;
    16'b0001000000000000: out_v[97] = 10'b0111110100;
    16'b0000000000000001: out_v[97] = 10'b0001111100;
    16'b1000010010000100: out_v[97] = 10'b1001001000;
    16'b1000000010000100: out_v[97] = 10'b1101001111;
    16'b0000000000100000: out_v[97] = 10'b1011100010;
    16'b0000010000100000: out_v[97] = 10'b1110000011;
    default: out_v[97] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0111010100110010: out_v[98] = 10'b1100001010;
    16'b0110000100000010: out_v[98] = 10'b0011111111;
    16'b0010010000010010: out_v[98] = 10'b1000011111;
    16'b0111010100000110: out_v[98] = 10'b1000011111;
    16'b0111010000100011: out_v[98] = 10'b0001110111;
    16'b0111010000110111: out_v[98] = 10'b0111100010;
    16'b0111010000010010: out_v[98] = 10'b1110111110;
    16'b0101000000000000: out_v[98] = 10'b1010011101;
    16'b0110010000010010: out_v[98] = 10'b1110110111;
    16'b0111010100000010: out_v[98] = 10'b1111110011;
    16'b0110010000110010: out_v[98] = 10'b1111101010;
    16'b0101010000110011: out_v[98] = 10'b0100100011;
    16'b0111000000000010: out_v[98] = 10'b1001000110;
    16'b0111010100110011: out_v[98] = 10'b1110001010;
    16'b0111010000110010: out_v[98] = 10'b1110101100;
    16'b0101010000110010: out_v[98] = 10'b0111001100;
    16'b0011010000110010: out_v[98] = 10'b1011011100;
    16'b0110010100010010: out_v[98] = 10'b0110110000;
    16'b0111010000110110: out_v[98] = 10'b0000010110;
    16'b0111010000110011: out_v[98] = 10'b0111001101;
    16'b0111010000000010: out_v[98] = 10'b1111010011;
    16'b1111000100000111: out_v[98] = 10'b1000101011;
    16'b0111010000101111: out_v[98] = 10'b0111111111;
    16'b0111000100000110: out_v[98] = 10'b1010111001;
    16'b0001010000110011: out_v[98] = 10'b1001111011;
    16'b0101000000010000: out_v[98] = 10'b1010011101;
    16'b0111000000000110: out_v[98] = 10'b1010011111;
    16'b0111000100000010: out_v[98] = 10'b0110001000;
    16'b0111010100100010: out_v[98] = 10'b1000110111;
    16'b0111000100000000: out_v[98] = 10'b0111110011;
    16'b0100000000000000: out_v[98] = 10'b0011110111;
    16'b0111010000100010: out_v[98] = 10'b1111010110;
    16'b0111010000100111: out_v[98] = 10'b1110101110;
    16'b0010010000110010: out_v[98] = 10'b1111011101;
    16'b0001010000110010: out_v[98] = 10'b0111110011;
    16'b0111010100010010: out_v[98] = 10'b1111011110;
    16'b0111000000000000: out_v[98] = 10'b0101101011;
    16'b0101010000110111: out_v[98] = 10'b1101110111;
    16'b0111010000000110: out_v[98] = 10'b1011000011;
    16'b1011000100000101: out_v[98] = 10'b0010011011;
    16'b0110010100110010: out_v[98] = 10'b0111001011;
    16'b0111010100110111: out_v[98] = 10'b1101110011;
    16'b1010000000000001: out_v[98] = 10'b0000111011;
    16'b0001000000000000: out_v[98] = 10'b1111101101;
    16'b0001000000000101: out_v[98] = 10'b1100000011;
    16'b0001000000000100: out_v[98] = 10'b0101001110;
    16'b0000000100000001: out_v[98] = 10'b1000010011;
    16'b0001000000000001: out_v[98] = 10'b0111010001;
    16'b0010000100000001: out_v[98] = 10'b1011100101;
    16'b0010000000000001: out_v[98] = 10'b1011001011;
    16'b0001000100000001: out_v[98] = 10'b0101001100;
    16'b0001000100000101: out_v[98] = 10'b1011011111;
    16'b0000000000000100: out_v[98] = 10'b1010001010;
    16'b0000000000000001: out_v[98] = 10'b0111110011;
    16'b1001000000000101: out_v[98] = 10'b0011110011;
    16'b0010000000000000: out_v[98] = 10'b1011011010;
    16'b1001000000000100: out_v[98] = 10'b1000001001;
    16'b1010000100000001: out_v[98] = 10'b0100001101;
    16'b1010000000000011: out_v[98] = 10'b0010110010;
    16'b0011000100000101: out_v[98] = 10'b1110111110;
    16'b0011000000000001: out_v[98] = 10'b0111011001;
    16'b0011000000000101: out_v[98] = 10'b0110010110;
    16'b1001000100000101: out_v[98] = 10'b0011101000;
    16'b0011000100000001: out_v[98] = 10'b1011010111;
    16'b1001000000000001: out_v[98] = 10'b1101001000;
    16'b1000000000000001: out_v[98] = 10'b0011101100;
    16'b1110000100010001: out_v[98] = 10'b0100111101;
    16'b1011000100000001: out_v[98] = 10'b0110011100;
    16'b0001000000010001: out_v[98] = 10'b0010110110;
    16'b0010000100000000: out_v[98] = 10'b1010000100;
    16'b1101000000010001: out_v[98] = 10'b1000100111;
    16'b1011000100000011: out_v[98] = 10'b0001111001;
    16'b1011000000000011: out_v[98] = 10'b1101000011;
    16'b1000000000000000: out_v[98] = 10'b0000011011;
    16'b1010000100100011: out_v[98] = 10'b1111101011;
    16'b1011000000000001: out_v[98] = 10'b0011101110;
    16'b1000000100000001: out_v[98] = 10'b0000111100;
    16'b1100000000010001: out_v[98] = 10'b1011001001;
    16'b1001000000010001: out_v[98] = 10'b0100111010;
    16'b1000000010000001: out_v[98] = 10'b1101001111;
    16'b1001000000000000: out_v[98] = 10'b1011000001;
    16'b1010000100000011: out_v[98] = 10'b1000100100;
    16'b1010000100010001: out_v[98] = 10'b1111101101;
    16'b1000000000010001: out_v[98] = 10'b0011100001;
    16'b0001000010000001: out_v[98] = 10'b1111111100;
    16'b0101000000010001: out_v[98] = 10'b0100010111;
    16'b1001100010000001: out_v[98] = 10'b0001001101;
    16'b1011000100100011: out_v[98] = 10'b1101010101;
    16'b0101000000010101: out_v[98] = 10'b1110010111;
    16'b1010000110000001: out_v[98] = 10'b0111111011;
    16'b1001000010000001: out_v[98] = 10'b0101111110;
    16'b1010000100000000: out_v[98] = 10'b1111000111;
    16'b1101000000000001: out_v[98] = 10'b1000101101;
    16'b1100000000000100: out_v[98] = 10'b1110100101;
    16'b1101000000000000: out_v[98] = 10'b1111010000;
    16'b1011000000000010: out_v[98] = 10'b1101001010;
    16'b1111000100000100: out_v[98] = 10'b1111001111;
    16'b1110000100000010: out_v[98] = 10'b1111110110;
    16'b1101000000000100: out_v[98] = 10'b1001001100;
    16'b1100000000000000: out_v[98] = 10'b0100101101;
    16'b1110000100000100: out_v[98] = 10'b1101011111;
    16'b1010000000000010: out_v[98] = 10'b1001011011;
    16'b1111000000000010: out_v[98] = 10'b1010001010;
    16'b1110000000000010: out_v[98] = 10'b1111000010;
    16'b1011000000000000: out_v[98] = 10'b1010001111;
    16'b1101000000010100: out_v[98] = 10'b1111000001;
    16'b1011000000000100: out_v[98] = 10'b0110110101;
    16'b0000000000000000: out_v[98] = 10'b0000011001;
    16'b1011000100000000: out_v[98] = 10'b0111000001;
    16'b1100000000010000: out_v[98] = 10'b1110111011;
    16'b1010000000000100: out_v[98] = 10'b0101011111;
    16'b1101000000010000: out_v[98] = 10'b0010011111;
    16'b1111000000000110: out_v[98] = 10'b0110100110;
    16'b1010000000000000: out_v[98] = 10'b0001111001;
    16'b0011000000000000: out_v[98] = 10'b0010100100;
    16'b1110000000000000: out_v[98] = 10'b0001010011;
    16'b1111000000000100: out_v[98] = 10'b0101100111;
    16'b1101000000010101: out_v[98] = 10'b1100011010;
    16'b0101000000000100: out_v[98] = 10'b1010011001;
    16'b0101000000010100: out_v[98] = 10'b0001011110;
    16'b1010000100000100: out_v[98] = 10'b0001011010;
    16'b1110000100000000: out_v[98] = 10'b1011011101;
    16'b1000000000000100: out_v[98] = 10'b1000101101;
    16'b1100000000010100: out_v[98] = 10'b1101100110;
    16'b1111000000000000: out_v[98] = 10'b0110110011;
    16'b1101000000000101: out_v[98] = 10'b1110001001;
    16'b1110000000000100: out_v[98] = 10'b0111100111;
    16'b1010000100000010: out_v[98] = 10'b1110010100;
    16'b1000000000001010: out_v[98] = 10'b1001100011;
    16'b1110000000000001: out_v[98] = 10'b1000000011;
    16'b1001000000000011: out_v[98] = 10'b1000011110;
    16'b1001000000001011: out_v[98] = 10'b0011011001;
    16'b1000000000000010: out_v[98] = 10'b0000011110;
    16'b1001000000001111: out_v[98] = 10'b0011110011;
    16'b1000000100000000: out_v[98] = 10'b0110110011;
    16'b1000000000000011: out_v[98] = 10'b1000101111;
    16'b1010000000100000: out_v[98] = 10'b0101101011;
    16'b1000000000001011: out_v[98] = 10'b0001111110;
    16'b1110000000100000: out_v[98] = 10'b0011101100;
    16'b1001000000000010: out_v[98] = 10'b0000111101;
    16'b1000000000101011: out_v[98] = 10'b1110010000;
    16'b1110000000100010: out_v[98] = 10'b0111101011;
    16'b1000000000101010: out_v[98] = 10'b0011111011;
    16'b1100000000000010: out_v[98] = 10'b0010101111;
    16'b1100000000101010: out_v[98] = 10'b1101001111;
    16'b0000000000000111: out_v[98] = 10'b1011101100;
    16'b0000000000001111: out_v[98] = 10'b0011100100;
    16'b1011000000001100: out_v[98] = 10'b1011010011;
    16'b0011000000001100: out_v[98] = 10'b1011010110;
    16'b0001000000001011: out_v[98] = 10'b1111011111;
    16'b1011000000001101: out_v[98] = 10'b1110100110;
    16'b0011000000001110: out_v[98] = 10'b1110110011;
    16'b1001000000000111: out_v[98] = 10'b0111111101;
    16'b0011000000001001: out_v[98] = 10'b1000111000;
    16'b0011000000001111: out_v[98] = 10'b1110110101;
    16'b0011000000001010: out_v[98] = 10'b1101010101;
    16'b1111000000010000: out_v[98] = 10'b0001110101;
    16'b0011000000001101: out_v[98] = 10'b0010111001;
    16'b1011000000001000: out_v[98] = 10'b0001011010;
    16'b0011000000001000: out_v[98] = 10'b0011011010;
    16'b1011000100000100: out_v[98] = 10'b1110110001;
    16'b0001000000001110: out_v[98] = 10'b1111001011;
    16'b0001000000001010: out_v[98] = 10'b1100000110;
    16'b1111000000001000: out_v[98] = 10'b1110110111;
    16'b0001000000001111: out_v[98] = 10'b1001111110;
    16'b0001000000000010: out_v[98] = 10'b0001100010;
    16'b0011000000000100: out_v[98] = 10'b1100100101;
    16'b1100000100000000: out_v[98] = 10'b0010101011;
    16'b0000000000000011: out_v[98] = 10'b1101101001;
    16'b0001000000000110: out_v[98] = 10'b1011100110;
    16'b1001000000001010: out_v[98] = 10'b0110011111;
    16'b0001000000000011: out_v[98] = 10'b1111111100;
    16'b0001000000000111: out_v[98] = 10'b1101111010;
    16'b1011000000001110: out_v[98] = 10'b1110010010;
    16'b1101000100010001: out_v[98] = 10'b1100110001;
    16'b1101000100000101: out_v[98] = 10'b0011100010;
    16'b1111000100010101: out_v[98] = 10'b1110110100;
    16'b1101000100000001: out_v[98] = 10'b1100001011;
    16'b1100010000010001: out_v[98] = 10'b1011001110;
    16'b1001000100000001: out_v[98] = 10'b1101110010;
    16'b1100000000000001: out_v[98] = 10'b1011101011;
    16'b1111000100000101: out_v[98] = 10'b1010111000;
    16'b1111000100000001: out_v[98] = 10'b0111011001;
    16'b1000010000010001: out_v[98] = 10'b0110111011;
    16'b1101000100010101: out_v[98] = 10'b1111010010;
    16'b0101000100000101: out_v[98] = 10'b0011100111;
    16'b1100010000000001: out_v[98] = 10'b1011101110;
    16'b1100000100010001: out_v[98] = 10'b0110111010;
    16'b1011000000000101: out_v[98] = 10'b1100110100;
    16'b1001000100000100: out_v[98] = 10'b1101011110;
    16'b1101010100010001: out_v[98] = 10'b1011110010;
    16'b1101000100000000: out_v[98] = 10'b1011110010;
    16'b0000010000010001: out_v[98] = 10'b1111010000;
    16'b0100000000000001: out_v[98] = 10'b1001000101;
    16'b1101000100000100: out_v[98] = 10'b1011011111;
    16'b1100000100000001: out_v[98] = 10'b1000111010;
    16'b0100010000010001: out_v[98] = 10'b1111101110;
    16'b1111000000000101: out_v[98] = 10'b0011111010;
    16'b0100000000010001: out_v[98] = 10'b1001010110;
    16'b1000000000000110: out_v[98] = 10'b1011101001;
    16'b1101000000000010: out_v[98] = 10'b0011100111;
    16'b1000000000000111: out_v[98] = 10'b0111001001;
    16'b1001000000000110: out_v[98] = 10'b0001111010;
    16'b1001001000000011: out_v[98] = 10'b1101110111;
    16'b1011000000001111: out_v[98] = 10'b0001110101;
    16'b1011000000000110: out_v[98] = 10'b0100101110;
    16'b1011000000000111: out_v[98] = 10'b1001000100;
    16'b1011000000001011: out_v[98] = 10'b1101001100;
    16'b1011000000001010: out_v[98] = 10'b0011010111;
    16'b1011010000000011: out_v[98] = 10'b1001101010;
    16'b0011000000000010: out_v[98] = 10'b0111011101;
    16'b0011000000000011: out_v[98] = 10'b0101011111;
    16'b1010000000000101: out_v[98] = 10'b0111001011;
    16'b0011000000000110: out_v[98] = 10'b1111010111;
    16'b1011000100000111: out_v[98] = 10'b1101110001;
    16'b1000000000000101: out_v[98] = 10'b0110100001;
    16'b1101100001000000: out_v[98] = 10'b1101010101;
    16'b1011000000100010: out_v[98] = 10'b1011101101;
    16'b1001000001000000: out_v[98] = 10'b1111001011;
    default: out_v[98] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1000111000000001: out_v[99] = 10'b0111111011;
    16'b0100110010010010: out_v[99] = 10'b1111111111;
    16'b0000110010000011: out_v[99] = 10'b1111110010;
    16'b0100110010000000: out_v[99] = 10'b1001001110;
    16'b0100111000000001: out_v[99] = 10'b1010110111;
    16'b0000011010000011: out_v[99] = 10'b0111100010;
    16'b0100100010000000: out_v[99] = 10'b0110110111;
    16'b1000101000000001: out_v[99] = 10'b0011010011;
    16'b0100110010000011: out_v[99] = 10'b1110111111;
    16'b0100111010000011: out_v[99] = 10'b1001011110;
    16'b1100110010000000: out_v[99] = 10'b1001001001;
    16'b0000100000000000: out_v[99] = 10'b0011000101;
    16'b0000101000000001: out_v[99] = 10'b0000101101;
    16'b1000100000000001: out_v[99] = 10'b0111110011;
    16'b1000001000000001: out_v[99] = 10'b1000011111;
    16'b0100110010000001: out_v[99] = 10'b1111101010;
    16'b0000111000000001: out_v[99] = 10'b1101110110;
    16'b1100111010000001: out_v[99] = 10'b1110001010;
    16'b0000110000000001: out_v[99] = 10'b1000101011;
    16'b0100110010010000: out_v[99] = 10'b0001100111;
    16'b1000111010000001: out_v[99] = 10'b1111000000;
    16'b0100010010000000: out_v[99] = 10'b0011101110;
    16'b0100111010000001: out_v[99] = 10'b0000110111;
    16'b0000110010000001: out_v[99] = 10'b0110110110;
    16'b0100100010000001: out_v[99] = 10'b1001000011;
    16'b0000110010000000: out_v[99] = 10'b1001101110;
    16'b0000100010000000: out_v[99] = 10'b1001110111;
    16'b0100110010000010: out_v[99] = 10'b1111011011;
    16'b0100010010000011: out_v[99] = 10'b1111111000;
    16'b0000111010000001: out_v[99] = 10'b1010010010;
    16'b0000110000000000: out_v[99] = 10'b0100111100;
    16'b0100010010000010: out_v[99] = 10'b1000111111;
    16'b1000110010000000: out_v[99] = 10'b1011111110;
    16'b0000110010000010: out_v[99] = 10'b1101110111;
    16'b0100010010000001: out_v[99] = 10'b0110111011;
    16'b0100011010000011: out_v[99] = 10'b1010110100;
    16'b0000111010000011: out_v[99] = 10'b1100111110;
    16'b1000100000000000: out_v[99] = 10'b0110000110;
    16'b1000110010000001: out_v[99] = 10'b1111111010;
    16'b0000101000000011: out_v[99] = 10'b1000110101;
    16'b0000001000000001: out_v[99] = 10'b0101001011;
    16'b0000100000000001: out_v[99] = 10'b1111000101;
    16'b0100110000000000: out_v[99] = 10'b1010010111;
    16'b1100111000000001: out_v[99] = 10'b1001000011;
    16'b1100110010000001: out_v[99] = 10'b1011111011;
    16'b0100100010000010: out_v[99] = 10'b0011100000;
    16'b0100110000000001: out_v[99] = 10'b0000110101;
    16'b0100001001000011: out_v[99] = 10'b0111011000;
    16'b0000000001000010: out_v[99] = 10'b1000000011;
    16'b1000000001000010: out_v[99] = 10'b0111010011;
    16'b0100001001010011: out_v[99] = 10'b0000110111;
    16'b0100011001000011: out_v[99] = 10'b0011110101;
    16'b0000000001000011: out_v[99] = 10'b1110101101;
    16'b0000100001000010: out_v[99] = 10'b0000011111;
    16'b1000100001000010: out_v[99] = 10'b0100011011;
    16'b0100001001000001: out_v[99] = 10'b0101001001;
    16'b0100011011000011: out_v[99] = 10'b1010011011;
    16'b0000001001000011: out_v[99] = 10'b1110001100;
    16'b0100000001000010: out_v[99] = 10'b0010100011;
    16'b0100000001000011: out_v[99] = 10'b0011001111;
    16'b0100011001010011: out_v[99] = 10'b0101000111;
    16'b0100000001000001: out_v[99] = 10'b1001011010;
    16'b0100000001000000: out_v[99] = 10'b0000111011;
    16'b1000101001000011: out_v[99] = 10'b0100111110;
    16'b0000101001000011: out_v[99] = 10'b0111000010;
    16'b0000101001000001: out_v[99] = 10'b1010011011;
    16'b0100101011000001: out_v[99] = 10'b0100101010;
    16'b0100101011000011: out_v[99] = 10'b1010111101;
    16'b0000001001000001: out_v[99] = 10'b1111000100;
    16'b0000100010000001: out_v[99] = 10'b1111010111;
    16'b0100011010000001: out_v[99] = 10'b0010000111;
    16'b0000000000000001: out_v[99] = 10'b1101000100;
    16'b0100111011000001: out_v[99] = 10'b1110110111;
    16'b0000000000000000: out_v[99] = 10'b0010010010;
    16'b0000000010000001: out_v[99] = 10'b0001100110;
    16'b0000101010000001: out_v[99] = 10'b1100010110;
    16'b0000001011000001: out_v[99] = 10'b1001100111;
    16'b0000101011000011: out_v[99] = 10'b0011001010;
    16'b0000001010000001: out_v[99] = 10'b0001011110;
    16'b0100111011000011: out_v[99] = 10'b1110111010;
    16'b0000101011000001: out_v[99] = 10'b0111010000;
    16'b0000000010000000: out_v[99] = 10'b1101101100;
    16'b0100101010000001: out_v[99] = 10'b0011110111;
    16'b0000101001000010: out_v[99] = 10'b0011010101;
    16'b0000001000000000: out_v[99] = 10'b1001001111;
    16'b0000100001000000: out_v[99] = 10'b1100001111;
    16'b0000001001000010: out_v[99] = 10'b1000101101;
    16'b0000001011000011: out_v[99] = 10'b1011100110;
    16'b0100101000000001: out_v[99] = 10'b0010011100;
    16'b1000101001000001: out_v[99] = 10'b0111101010;
    16'b0100000010000001: out_v[99] = 10'b1011011011;
    16'b0100001010000001: out_v[99] = 10'b1100000111;
    16'b1000000000000000: out_v[99] = 10'b0100010111;
    16'b0100011011000001: out_v[99] = 10'b1011111111;
    16'b0100101001000011: out_v[99] = 10'b0001110110;
    16'b0000000001000000: out_v[99] = 10'b1001011001;
    16'b1000000001000000: out_v[99] = 10'b1100101010;
    16'b0100110001000010: out_v[99] = 10'b1100001011;
    16'b1000100001010010: out_v[99] = 10'b0011011111;
    16'b0100110001010010: out_v[99] = 10'b0001011011;
    16'b0100110011000010: out_v[99] = 10'b0011001111;
    16'b1000100000000010: out_v[99] = 10'b0010111000;
    16'b1000100001000011: out_v[99] = 10'b1011011001;
    16'b0000100011000010: out_v[99] = 10'b0110001011;
    16'b1000100011000010: out_v[99] = 10'b0000011101;
    16'b0100110011000000: out_v[99] = 10'b1011101110;
    16'b0000110001010010: out_v[99] = 10'b0101100111;
    16'b1100110011000010: out_v[99] = 10'b0110010111;
    16'b0000000001010010: out_v[99] = 10'b0101100110;
    16'b0100010001010010: out_v[99] = 10'b0111010010;
    16'b0100000011000010: out_v[99] = 10'b1111111000;
    16'b0000100011000011: out_v[99] = 10'b1111011011;
    16'b0100010011000011: out_v[99] = 10'b0110011001;
    16'b0100100011000010: out_v[99] = 10'b0110110111;
    16'b0100110011000011: out_v[99] = 10'b1001011101;
    16'b1000100001000000: out_v[99] = 10'b1100100001;
    16'b0000100001010010: out_v[99] = 10'b0111011111;
    16'b0000100000000010: out_v[99] = 10'b0011111100;
    16'b0100010011000010: out_v[99] = 10'b0110010101;
    16'b0100100001000010: out_v[99] = 10'b0101100100;
    16'b0100100011000011: out_v[99] = 10'b1011000011;
    16'b1000100011000011: out_v[99] = 10'b1011001111;
    16'b0100110011010010: out_v[99] = 10'b1011001011;
    16'b1100100011000010: out_v[99] = 10'b0011111111;
    16'b0000100001000011: out_v[99] = 10'b0100001011;
    16'b0000000000000010: out_v[99] = 10'b1010100000;
    16'b0000010001000010: out_v[99] = 10'b1001010101;
    16'b0100010000000000: out_v[99] = 10'b1010011010;
    16'b0000010001000000: out_v[99] = 10'b1100000111;
    16'b0001010000000000: out_v[99] = 10'b0011011100;
    16'b0100000000000000: out_v[99] = 10'b0010110011;
    16'b0000010000000000: out_v[99] = 10'b0011110010;
    16'b1100000000000000: out_v[99] = 10'b1000111101;
    16'b0100100000000000: out_v[99] = 10'b0000110101;
    16'b1000110000000000: out_v[99] = 10'b0110110110;
    16'b1100100000000000: out_v[99] = 10'b0001110110;
    16'b1100110001000000: out_v[99] = 10'b1111111101;
    16'b1000010000000000: out_v[99] = 10'b1010001001;
    16'b1100110000000000: out_v[99] = 10'b0111011010;
    16'b1100100001000000: out_v[99] = 10'b1011100011;
    16'b1000110001000000: out_v[99] = 10'b1111110010;
    16'b0001000000000000: out_v[99] = 10'b0001111011;
    16'b0100010001000000: out_v[99] = 10'b1101101110;
    16'b0001010001000000: out_v[99] = 10'b1111000111;
    16'b0100000000000010: out_v[99] = 10'b0000110101;
    16'b0000010000000010: out_v[99] = 10'b1110001000;
    16'b0001000001000000: out_v[99] = 10'b0101010111;
    16'b1100100001000010: out_v[99] = 10'b1110010001;
    16'b0001010011000011: out_v[99] = 10'b1011001111;
    16'b0001010011000010: out_v[99] = 10'b1011001111;
    16'b0000010011000011: out_v[99] = 10'b0100110011;
    16'b0100100001000000: out_v[99] = 10'b1110110010;
    16'b0100100011000000: out_v[99] = 10'b1111011000;
    16'b0000011011000011: out_v[99] = 10'b0010011001;
    16'b1100100001000011: out_v[99] = 10'b0100100110;
    16'b1100100001000001: out_v[99] = 10'b1000111111;
    16'b0000010010000011: out_v[99] = 10'b0000111011;
    16'b1100000001000000: out_v[99] = 10'b0010100101;
    16'b0100101000000011: out_v[99] = 10'b0111110010;
    16'b0100001000000011: out_v[99] = 10'b0001000001;
    16'b0000101000000000: out_v[99] = 10'b1100000101;
    16'b0100101001000001: out_v[99] = 10'b1111110010;
    16'b0000101001000000: out_v[99] = 10'b0001101101;
    16'b0000001001000000: out_v[99] = 10'b1001110011;
    16'b0000101000000010: out_v[99] = 10'b0001001011;
    16'b0000001000000011: out_v[99] = 10'b0000001111;
    16'b0000010000010010: out_v[99] = 10'b0010010101;
    16'b1000000000000010: out_v[99] = 10'b1000111000;
    16'b0000010000010000: out_v[99] = 10'b0111010011;
    16'b0000011001010001: out_v[99] = 10'b1110100011;
    16'b0000010000010001: out_v[99] = 10'b0111100111;
    16'b0000011000010001: out_v[99] = 10'b0101110011;
    16'b0000010000010011: out_v[99] = 10'b0110011100;
    16'b1000110000000010: out_v[99] = 10'b0001101101;
    16'b0000000000010000: out_v[99] = 10'b1011001010;
    16'b1000001001000001: out_v[99] = 10'b0101010100;
    16'b1000111001000001: out_v[99] = 10'b0011110101;
    16'b0100111001000001: out_v[99] = 10'b1011110110;
    16'b0000011001000011: out_v[99] = 10'b0101000101;
    16'b0100010011010010: out_v[99] = 10'b1111010101;
    16'b1100111001000001: out_v[99] = 10'b1101001000;
    16'b0000011001000001: out_v[99] = 10'b1100111011;
    16'b1100111001000011: out_v[99] = 10'b1001110101;
    16'b0100011001000001: out_v[99] = 10'b0111111010;
    16'b1000111001000011: out_v[99] = 10'b1100011011;
    16'b0100011000000001: out_v[99] = 10'b1000011011;
    16'b1100101001000011: out_v[99] = 10'b1110111011;
    16'b1000110001000010: out_v[99] = 10'b1100100100;
    16'b0100111001000011: out_v[99] = 10'b0010111001;
    16'b0100010001000010: out_v[99] = 10'b1101001100;
    16'b1000001001000011: out_v[99] = 10'b0111110010;
    16'b1100101001000001: out_v[99] = 10'b0111011011;
    16'b1000101000000000: out_v[99] = 10'b1100001011;
    16'b0000010001010001: out_v[99] = 10'b0111100111;
    16'b0000010001010000: out_v[99] = 10'b1001011011;
    default: out_v[99] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010000010000000: out_v[100] = 10'b1111011010;
    16'b1010000110010000: out_v[100] = 10'b1011000001;
    16'b1010001110110000: out_v[100] = 10'b1100010011;
    16'b1010001010110000: out_v[100] = 10'b1111001110;
    16'b1010000010100000: out_v[100] = 10'b0111000011;
    16'b1000001010100000: out_v[100] = 10'b1100011001;
    16'b0010001110010000: out_v[100] = 10'b0011111011;
    16'b1010001110010000: out_v[100] = 10'b1101011101;
    16'b1010000010010000: out_v[100] = 10'b0111001101;
    16'b1010001100000000: out_v[100] = 10'b0010000101;
    16'b1010000010000000: out_v[100] = 10'b1011010011;
    16'b1010000010110000: out_v[100] = 10'b1010110000;
    16'b1010000110110000: out_v[100] = 10'b0111011010;
    16'b1010001010100000: out_v[100] = 10'b0111000100;
    16'b0010000010010000: out_v[100] = 10'b1000111011;
    16'b0010000100010000: out_v[100] = 10'b1100001011;
    16'b1010001110100000: out_v[100] = 10'b1010100100;
    16'b1000001110110000: out_v[100] = 10'b1001011111;
    16'b0010000110010000: out_v[100] = 10'b1100000100;
    16'b1000001010110000: out_v[100] = 10'b0001001011;
    16'b0000000010010000: out_v[100] = 10'b1100000100;
    16'b1010001010010000: out_v[100] = 10'b1011000111;
    16'b0010000010100000: out_v[100] = 10'b1100000001;
    16'b0010000000010000: out_v[100] = 10'b1011111001;
    16'b0000000010000000: out_v[100] = 10'b1100100001;
    16'b1000001110100000: out_v[100] = 10'b0101110111;
    16'b0000000000010000: out_v[100] = 10'b0110100011;
    16'b0000000000000000: out_v[100] = 10'b0111001111;
    16'b0000000010000100: out_v[100] = 10'b1111011101;
    16'b0000000010010100: out_v[100] = 10'b0110110110;
    16'b1000000010010000: out_v[100] = 10'b1011100010;
    16'b1000000000010001: out_v[100] = 10'b1110010011;
    16'b0000000000010001: out_v[100] = 10'b1011111000;
    16'b1000000010010100: out_v[100] = 10'b1111011011;
    16'b1000000010000000: out_v[100] = 10'b1010110100;
    16'b1000000000100000: out_v[100] = 10'b1000001101;
    16'b0000000010010001: out_v[100] = 10'b0000011001;
    16'b0010001000000000: out_v[100] = 10'b0011010101;
    16'b1000000000000000: out_v[100] = 10'b1101000110;
    16'b1100000000000100: out_v[100] = 10'b0111001001;
    16'b0000000000110000: out_v[100] = 10'b0011011001;
    16'b1000000010110000: out_v[100] = 10'b0011101100;
    16'b1100000010000100: out_v[100] = 10'b1100101110;
    16'b0000000000000001: out_v[100] = 10'b1110110101;
    16'b1000000000010000: out_v[100] = 10'b1010000111;
    16'b1000000000000100: out_v[100] = 10'b1010101000;
    16'b1010001000000000: out_v[100] = 10'b1001100111;
    16'b1100000000010100: out_v[100] = 10'b1001001110;
    16'b0100000010000100: out_v[100] = 10'b0110110111;
    16'b0000000010100000: out_v[100] = 10'b0110101100;
    16'b1100000000000000: out_v[100] = 10'b1001101001;
    16'b1100000010010100: out_v[100] = 10'b0000001010;
    16'b0010000000000000: out_v[100] = 10'b0010110011;
    16'b0000000010110000: out_v[100] = 10'b1000110110;
    16'b1000000010100000: out_v[100] = 10'b0000001101;
    16'b1000000000000001: out_v[100] = 10'b0010110001;
    16'b0100000010010100: out_v[100] = 10'b0100000110;
    16'b1000000000010100: out_v[100] = 10'b1100011101;
    16'b0100000000000100: out_v[100] = 10'b0110000101;
    16'b1000000000110000: out_v[100] = 10'b1000001101;
    16'b0000000000000100: out_v[100] = 10'b0000110011;
    16'b1000000010000100: out_v[100] = 10'b1001011010;
    16'b0000000010000001: out_v[100] = 10'b1001001100;
    16'b1000000010000001: out_v[100] = 10'b1101100010;
    16'b1000000010010001: out_v[100] = 10'b0111100101;
    16'b1010000000000000: out_v[100] = 10'b1000011011;
    16'b0000000000100000: out_v[100] = 10'b0110001100;
    16'b0010000010010100: out_v[100] = 10'b0111011110;
    16'b1110000010010100: out_v[100] = 10'b0001001101;
    16'b1100000010010000: out_v[100] = 10'b0011111010;
    16'b1010000010010100: out_v[100] = 10'b0011001011;
    16'b1110000010010000: out_v[100] = 10'b1111011011;
    16'b1110000010000100: out_v[100] = 10'b1001001010;
    16'b1110000010000000: out_v[100] = 10'b1111010100;
    16'b1100000010000000: out_v[100] = 10'b1000011100;
    16'b0100000000000000: out_v[100] = 10'b1101001111;
    16'b1010000010000100: out_v[100] = 10'b1010011000;
    16'b0010000000100000: out_v[100] = 10'b1001010101;
    16'b0010001010000000: out_v[100] = 10'b0010111100;
    16'b0010001000100000: out_v[100] = 10'b0111111011;
    16'b0110000000000000: out_v[100] = 10'b1001110011;
    16'b0010001010100000: out_v[100] = 10'b0001111000;
    16'b0000001010100000: out_v[100] = 10'b0100110011;
    16'b1010000000100000: out_v[100] = 10'b1110100000;
    16'b1010001000100000: out_v[100] = 10'b0100001010;
    16'b1100001000000000: out_v[100] = 10'b1111110000;
    16'b0000001000100000: out_v[100] = 10'b1101100011;
    16'b1110001000000000: out_v[100] = 10'b1001111010;
    16'b0010001110000000: out_v[100] = 10'b0100010110;
    16'b0010000000100100: out_v[100] = 10'b1101011010;
    16'b0000001000000000: out_v[100] = 10'b1100010010;
    16'b0110001000000000: out_v[100] = 10'b0011111010;
    16'b1000001000100000: out_v[100] = 10'b1010100010;
    16'b0010100000000000: out_v[100] = 10'b0111100110;
    16'b0010000010110000: out_v[100] = 10'b0111110001;
    16'b0000000100000000: out_v[100] = 10'b0010111010;
    16'b0010100010000000: out_v[100] = 10'b1000100110;
    16'b0010100010010000: out_v[100] = 10'b1011111110;
    16'b0010100010110000: out_v[100] = 10'b1111010111;
    16'b0010000100000000: out_v[100] = 10'b1000101001;
    16'b1010000010100100: out_v[100] = 10'b0011110011;
    16'b1010000010110100: out_v[100] = 10'b0010100111;
    16'b0010100010100000: out_v[100] = 10'b0010101111;
    16'b0010000110000000: out_v[100] = 10'b0100110000;
    16'b0000100010010000: out_v[100] = 10'b1100010110;
    16'b0010000000000001: out_v[100] = 10'b1101100010;
    16'b1010000000100010: out_v[100] = 10'b1111100010;
    16'b1010000000100001: out_v[100] = 10'b1010101001;
    16'b1010000010000001: out_v[100] = 10'b1011010110;
    16'b1010000000100110: out_v[100] = 10'b1111111001;
    16'b0010000010000001: out_v[100] = 10'b0111000111;
    16'b1010001000100001: out_v[100] = 10'b1000011011;
    16'b1010000010100001: out_v[100] = 10'b0101011110;
    16'b1010000000000001: out_v[100] = 10'b1111100111;
    16'b0100000010000000: out_v[100] = 10'b0110100010;
    16'b0000000110100000: out_v[100] = 10'b0011101011;
    16'b1100000000100000: out_v[100] = 10'b0010101111;
    16'b0100000010100000: out_v[100] = 10'b1010010100;
    16'b0100000000100000: out_v[100] = 10'b0000001010;
    16'b1100000010100000: out_v[100] = 10'b1011000000;
    16'b0010000110100000: out_v[100] = 10'b1100011111;
    16'b0000000110010000: out_v[100] = 10'b1100000010;
    16'b0000000110000000: out_v[100] = 10'b0110111111;
    16'b0010000110110000: out_v[100] = 10'b0110101010;
    16'b0000000110110000: out_v[100] = 10'b1011011111;
    16'b0000000100010000: out_v[100] = 10'b1101110010;
    default: out_v[100] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000100110000: out_v[101] = 10'b1100001011;
    16'b0000000100100000: out_v[101] = 10'b0100010101;
    16'b1000000100100000: out_v[101] = 10'b0001111011;
    16'b0000000000110000: out_v[101] = 10'b0011101110;
    16'b1000000000110000: out_v[101] = 10'b0100000001;
    16'b1000000000100000: out_v[101] = 10'b0100001110;
    16'b0000000100000000: out_v[101] = 10'b1010010111;
    16'b0000000000100000: out_v[101] = 10'b0010100111;
    16'b0000000100010000: out_v[101] = 10'b1000111111;
    16'b0000000000000000: out_v[101] = 10'b0010101010;
    16'b1000000100110000: out_v[101] = 10'b1001110101;
    16'b0000000110100000: out_v[101] = 10'b0111010001;
    16'b0001000100100000: out_v[101] = 10'b0101000011;
    16'b1000000000010000: out_v[101] = 10'b0000010110;
    16'b0000000000010000: out_v[101] = 10'b0100111110;
    16'b0000000010000000: out_v[101] = 10'b0101001001;
    16'b1000000000000000: out_v[101] = 10'b0010011000;
    16'b0000000000100001: out_v[101] = 10'b0011011101;
    16'b1001000000100000: out_v[101] = 10'b0110110110;
    16'b1000000000100001: out_v[101] = 10'b1011111100;
    16'b1001000000110000: out_v[101] = 10'b1100011101;
    16'b1000000000111000: out_v[101] = 10'b0101011010;
    16'b1000000000110001: out_v[101] = 10'b1001011100;
    16'b0001000000100000: out_v[101] = 10'b0000111111;
    16'b1001000000000000: out_v[101] = 10'b0110100110;
    16'b0000000000110001: out_v[101] = 10'b1010100110;
    16'b1000000010100000: out_v[101] = 10'b0000001101;
    16'b1000000000011000: out_v[101] = 10'b0101100111;
    16'b0000000010110000: out_v[101] = 10'b1111010100;
    16'b1000000010110000: out_v[101] = 10'b1111001010;
    16'b1000000010010000: out_v[101] = 10'b1001010000;
    16'b1000000000101000: out_v[101] = 10'b1010001000;
    16'b1001000000010000: out_v[101] = 10'b0010011001;
    16'b1000001000100000: out_v[101] = 10'b1011100111;
    16'b1000000010000000: out_v[101] = 10'b1110000001;
    16'b0000000010010000: out_v[101] = 10'b0011110010;
    16'b0000000010100000: out_v[101] = 10'b1010100110;
    16'b1000000100010000: out_v[101] = 10'b0011110000;
    16'b1001000100010000: out_v[101] = 10'b1011011011;
    16'b1000000100000000: out_v[101] = 10'b0011100000;
    16'b1000000110010000: out_v[101] = 10'b0110111110;
    16'b0000000000110010: out_v[101] = 10'b1011001000;
    16'b1000000100010001: out_v[101] = 10'b1011001010;
    16'b1000000100100001: out_v[101] = 10'b1011001010;
    16'b1000000000010001: out_v[101] = 10'b1011100111;
    16'b1000000100110001: out_v[101] = 10'b1111010100;
    16'b1001000010000000: out_v[101] = 10'b0010010010;
    16'b0001000000000000: out_v[101] = 10'b0101010101;
    default: out_v[101] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000001011000000: out_v[102] = 10'b1001101010;
    16'b0000000011000000: out_v[102] = 10'b0000000111;
    16'b0000011011001000: out_v[102] = 10'b1011100011;
    16'b0000011011000000: out_v[102] = 10'b0011001111;
    16'b0000011010000000: out_v[102] = 10'b0011111000;
    16'b0000001001000000: out_v[102] = 10'b1110010001;
    16'b0000010000000000: out_v[102] = 10'b0010001101;
    16'b0000000000000000: out_v[102] = 10'b0011110110;
    16'b0000000010000000: out_v[102] = 10'b0010110101;
    16'b0000001010000000: out_v[102] = 10'b0111101010;
    16'b0000001001001000: out_v[102] = 10'b0111110111;
    16'b0000011000000000: out_v[102] = 10'b0000110111;
    16'b0000010011000000: out_v[102] = 10'b0100110110;
    16'b0000010010000000: out_v[102] = 10'b1000011111;
    16'b0000000001001000: out_v[102] = 10'b1110100001;
    16'b0000000010001000: out_v[102] = 10'b1001001010;
    16'b0000001011001000: out_v[102] = 10'b1001010000;
    16'b0000000001000000: out_v[102] = 10'b1010100110;
    16'b0000000011001000: out_v[102] = 10'b0011001011;
    16'b0000001000000000: out_v[102] = 10'b1110101000;
    16'b0000011010001000: out_v[102] = 10'b1100111010;
    16'b0000011001000000: out_v[102] = 10'b0110010011;
    16'b0000000000001000: out_v[102] = 10'b1110001010;
    16'b1000000010001000: out_v[102] = 10'b0010110110;
    16'b0000010000001000: out_v[102] = 10'b1001010100;
    16'b0000000000010000: out_v[102] = 10'b0000000110;
    16'b0000010000010000: out_v[102] = 10'b1101010010;
    16'b0000010010001000: out_v[102] = 10'b1001001111;
    16'b0000010001000000: out_v[102] = 10'b1101110101;
    16'b1000000000001000: out_v[102] = 10'b1100010101;
    16'b0000010000011000: out_v[102] = 10'b0000110110;
    16'b1000010000000000: out_v[102] = 10'b0111101011;
    16'b1000000000000000: out_v[102] = 10'b1000010101;
    16'b0000000010010000: out_v[102] = 10'b0011000111;
    16'b0010000000001000: out_v[102] = 10'b1000100111;
    16'b1000000010000000: out_v[102] = 10'b1000010110;
    16'b0000000000011000: out_v[102] = 10'b1010101100;
    16'b0000000001010000: out_v[102] = 10'b1111100110;
    16'b0000010001001000: out_v[102] = 10'b0001011000;
    16'b0010010000001000: out_v[102] = 10'b0111100100;
    16'b0000011000001000: out_v[102] = 10'b1111000111;
    16'b0000010010011000: out_v[102] = 10'b1111110111;
    16'b0000000010011000: out_v[102] = 10'b0101101000;
    16'b0000010011001000: out_v[102] = 10'b1001001000;
    16'b0000001010001000: out_v[102] = 10'b1100100100;
    16'b0000001000001000: out_v[102] = 10'b1000110100;
    16'b1000010001000000: out_v[102] = 10'b0000011011;
    16'b0000011001001000: out_v[102] = 10'b0111000001;
    16'b0000000001011000: out_v[102] = 10'b1001001110;
    16'b0000011001010000: out_v[102] = 10'b1011011100;
    16'b0000000011011000: out_v[102] = 10'b1101000110;
    16'b0000011000010000: out_v[102] = 10'b1011101011;
    16'b0000010001010000: out_v[102] = 10'b1111010011;
    16'b0000001001011000: out_v[102] = 10'b0011110010;
    16'b0000001001010000: out_v[102] = 10'b0110111010;
    16'b0000001000010000: out_v[102] = 10'b1011101011;
    16'b0000011011010000: out_v[102] = 10'b1111011111;
    16'b0000000011010000: out_v[102] = 10'b1100011111;
    16'b0000011001011000: out_v[102] = 10'b1111000111;
    16'b0000000000000010: out_v[102] = 10'b0111000110;
    default: out_v[102] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100000000000000: out_v[103] = 10'b1011100000;
    16'b0100001000000001: out_v[103] = 10'b1110011100;
    16'b0000001000000001: out_v[103] = 10'b0100000010;
    16'b0000001000000000: out_v[103] = 10'b1101000011;
    16'b0100000000001000: out_v[103] = 10'b0110011010;
    16'b0010001000001001: out_v[103] = 10'b1001001011;
    16'b0000000000000001: out_v[103] = 10'b0000001001;
    16'b0100001000001001: out_v[103] = 10'b0000101101;
    16'b0100001000000000: out_v[103] = 10'b1100010101;
    16'b0000001000001001: out_v[103] = 10'b0001110011;
    16'b0000000000000000: out_v[103] = 10'b1101100110;
    16'b1000001000000001: out_v[103] = 10'b1010010011;
    16'b0000001000001000: out_v[103] = 10'b0100011010;
    16'b0000001010000001: out_v[103] = 10'b0110000111;
    16'b0000000000001000: out_v[103] = 10'b0100011100;
    16'b1010001000000001: out_v[103] = 10'b1010011011;
    16'b0010001000000001: out_v[103] = 10'b0011000011;
    16'b1000001010000001: out_v[103] = 10'b0011010011;
    16'b0100001000001000: out_v[103] = 10'b1011100011;
    16'b0000000010000000: out_v[103] = 10'b0001100110;
    16'b1100000000000000: out_v[103] = 10'b0001111000;
    16'b0010000000001000: out_v[103] = 10'b0000011110;
    16'b1010000000000000: out_v[103] = 10'b1110001101;
    16'b1100000000001000: out_v[103] = 10'b1111001000;
    16'b1100001000000001: out_v[103] = 10'b1100011110;
    16'b1000000000001000: out_v[103] = 10'b0101011100;
    16'b1010000000001000: out_v[103] = 10'b1110000100;
    16'b0110000000001000: out_v[103] = 10'b1000011110;
    16'b0010000000000000: out_v[103] = 10'b1110000100;
    16'b1110000000001000: out_v[103] = 10'b0111001100;
    16'b0000000010001000: out_v[103] = 10'b1001101100;
    16'b1100001000000000: out_v[103] = 10'b0011010111;
    16'b0110000000000000: out_v[103] = 10'b0011101010;
    16'b0100000010000000: out_v[103] = 10'b1010011000;
    16'b0100000010001000: out_v[103] = 10'b1011010010;
    16'b1100000010001000: out_v[103] = 10'b0010000010;
    16'b1100000010000000: out_v[103] = 10'b0011110011;
    16'b1000000010001000: out_v[103] = 10'b0100111111;
    16'b0100001010000000: out_v[103] = 10'b1100001110;
    16'b0100001010001000: out_v[103] = 10'b1001100011;
    16'b0100001010001001: out_v[103] = 10'b0101010000;
    16'b0100001010000001: out_v[103] = 10'b1101011010;
    16'b1000001000001001: out_v[103] = 10'b0111000110;
    16'b1100001000001001: out_v[103] = 10'b0010111010;
    16'b1100001010001000: out_v[103] = 10'b1001011011;
    16'b1100001000001000: out_v[103] = 10'b0110100111;
    default: out_v[103] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001010000000000: out_v[104] = 10'b1100011001;
    16'b0000000000000100: out_v[104] = 10'b1000110101;
    16'b0000010000100100: out_v[104] = 10'b0010100101;
    16'b0000010000100110: out_v[104] = 10'b0110111000;
    16'b0000010000000000: out_v[104] = 10'b1001000101;
    16'b0000010000100000: out_v[104] = 10'b0000001001;
    16'b0000000000100110: out_v[104] = 10'b0011010111;
    16'b0001010100000000: out_v[104] = 10'b1000110011;
    16'b0000010000110000: out_v[104] = 10'b0001110010;
    16'b0000010000100010: out_v[104] = 10'b0110100001;
    16'b0000010000100111: out_v[104] = 10'b1110101110;
    16'b0000000000100100: out_v[104] = 10'b0000011011;
    16'b0001010100000100: out_v[104] = 10'b0011000101;
    16'b0000010000000100: out_v[104] = 10'b0111101110;
    16'b0001010000000100: out_v[104] = 10'b0110011011;
    16'b0000000000100111: out_v[104] = 10'b1001100001;
    16'b0001010000000111: out_v[104] = 10'b1101110001;
    16'b0001000000000100: out_v[104] = 10'b0111100011;
    16'b0001010000100100: out_v[104] = 10'b0111111111;
    16'b0001010000100111: out_v[104] = 10'b1111101111;
    16'b0000010000110100: out_v[104] = 10'b0000110101;
    16'b0001010000100000: out_v[104] = 10'b1101100000;
    16'b0001010000010100: out_v[104] = 10'b0110000111;
    16'b0000011100010100: out_v[104] = 10'b1010010111;
    16'b0000001000010000: out_v[104] = 10'b0110001111;
    16'b0000011000010100: out_v[104] = 10'b1110010101;
    16'b0000011000010000: out_v[104] = 10'b0110000011;
    16'b0000001000000000: out_v[104] = 10'b0000100010;
    16'b0000011000010001: out_v[104] = 10'b0110110011;
    16'b0000001000010100: out_v[104] = 10'b0100101010;
    16'b0000011100010000: out_v[104] = 10'b0100010100;
    16'b0000001100010000: out_v[104] = 10'b0010010101;
    16'b0001011000000000: out_v[104] = 10'b0100101110;
    16'b0001011100000000: out_v[104] = 10'b1001101000;
    16'b0000011100000000: out_v[104] = 10'b0110001000;
    16'b0000010100000000: out_v[104] = 10'b1001010101;
    16'b0000001100000000: out_v[104] = 10'b1101001010;
    16'b0001011100010100: out_v[104] = 10'b1010110010;
    16'b0000011100000100: out_v[104] = 10'b0110010000;
    16'b0001011000000010: out_v[104] = 10'b1011101110;
    16'b0000011100010010: out_v[104] = 10'b1101010010;
    16'b0001011100100000: out_v[104] = 10'b0001000110;
    16'b0000011100000010: out_v[104] = 10'b0001011001;
    16'b0001011100000010: out_v[104] = 10'b0111001011;
    16'b0100011000010000: out_v[104] = 10'b1111000011;
    16'b0000011000000000: out_v[104] = 10'b1001101010;
    16'b0000010100000100: out_v[104] = 10'b0011010100;
    16'b0001011100010000: out_v[104] = 10'b1101101100;
    16'b0001001000000100: out_v[104] = 10'b1000100110;
    16'b0000011100000011: out_v[104] = 10'b1010111111;
    16'b0001011100000011: out_v[104] = 10'b1111111011;
    16'b0001010000000011: out_v[104] = 10'b1011111101;
    16'b0000010000010000: out_v[104] = 10'b0111110110;
    16'b0001011000000011: out_v[104] = 10'b1011011101;
    16'b0001011000000100: out_v[104] = 10'b1101010110;
    16'b0000011100010011: out_v[104] = 10'b1011110111;
    16'b0100011100010000: out_v[104] = 10'b1111110100;
    16'b0001011100000100: out_v[104] = 10'b1100110110;
    16'b0001010000000010: out_v[104] = 10'b0110101111;
    16'b0001011100110000: out_v[104] = 10'b1101111010;
    16'b0000011000110000: out_v[104] = 10'b1001000100;
    16'b0001011100000111: out_v[104] = 10'b1001111011;
    16'b0001000100010101: out_v[104] = 10'b1111100110;
    16'b0001010100010111: out_v[104] = 10'b0111011111;
    16'b0001000000010100: out_v[104] = 10'b1111101111;
    16'b0001000100010111: out_v[104] = 10'b1110110111;
    16'b0001000100010000: out_v[104] = 10'b1110110110;
    16'b0001010100010100: out_v[104] = 10'b1010101111;
    16'b0000001100010100: out_v[104] = 10'b1101001010;
    16'b0000000100110100: out_v[104] = 10'b0101011000;
    16'b0001000100010100: out_v[104] = 10'b1100110010;
    16'b0001000100010110: out_v[104] = 10'b0111011111;
    16'b0001011000010000: out_v[104] = 10'b0011000100;
    16'b0001000000010000: out_v[104] = 10'b1001101011;
    16'b0001001000010100: out_v[104] = 10'b1101000011;
    16'b0001011000010100: out_v[104] = 10'b0111011011;
    16'b0001011100010111: out_v[104] = 10'b1011111111;
    16'b0001001100010100: out_v[104] = 10'b0011001010;
    16'b0001011100010010: out_v[104] = 10'b1011001010;
    16'b0000010100110000: out_v[104] = 10'b0000111010;
    16'b0001001100010111: out_v[104] = 10'b0110001010;
    16'b1001000100010101: out_v[104] = 10'b1011101011;
    16'b0001010100010000: out_v[104] = 10'b0110101001;
    16'b0000010100010100: out_v[104] = 10'b1000001101;
    16'b0000000000010100: out_v[104] = 10'b0000111010;
    16'b0001001100010101: out_v[104] = 10'b0011011111;
    16'b0001001000010000: out_v[104] = 10'b0110111001;
    16'b0001010100010110: out_v[104] = 10'b1111100110;
    16'b0000000100010100: out_v[104] = 10'b1001100101;
    16'b0000000000010000: out_v[104] = 10'b1001110100;
    16'b0001010100010010: out_v[104] = 10'b1110101110;
    16'b0001010000010000: out_v[104] = 10'b0101001001;
    16'b0000001000010101: out_v[104] = 10'b0101011001;
    16'b0000001000000100: out_v[104] = 10'b0001100110;
    16'b0000010100010000: out_v[104] = 10'b1101111010;
    16'b0001001100010000: out_v[104] = 10'b1011010111;
    16'b0000010000010100: out_v[104] = 10'b0111101100;
    16'b0001001100000000: out_v[104] = 10'b1001001111;
    16'b0001001100110000: out_v[104] = 10'b0010100010;
    16'b0001001000100000: out_v[104] = 10'b1011011111;
    16'b0000000100010000: out_v[104] = 10'b1101001011;
    16'b0001001000000000: out_v[104] = 10'b1000010000;
    16'b0000000100000000: out_v[104] = 10'b0010010010;
    16'b0001001100100000: out_v[104] = 10'b0110010110;
    16'b0001001100000100: out_v[104] = 10'b1001100110;
    16'b0000001100000100: out_v[104] = 10'b1101001000;
    16'b0001001000110000: out_v[104] = 10'b0010001001;
    16'b0001000000000000: out_v[104] = 10'b1111000010;
    16'b0001000100000000: out_v[104] = 10'b0011010001;
    16'b0001000100100000: out_v[104] = 10'b0100111010;
    16'b0000001000000101: out_v[104] = 10'b1111111111;
    16'b0000000000000000: out_v[104] = 10'b1101100000;
    16'b0000011000000100: out_v[104] = 10'b1000110110;
    16'b0000011000000010: out_v[104] = 10'b1100011001;
    16'b0000011000010010: out_v[104] = 10'b1100110111;
    16'b0000000000110100: out_v[104] = 10'b0001110111;
    16'b0000010100110100: out_v[104] = 10'b1111001110;
    16'b0001011000100000: out_v[104] = 10'b0100100100;
    16'b0000011100100000: out_v[104] = 10'b0101101010;
    16'b0000011100110000: out_v[104] = 10'b1101001010;
    16'b0001010100100000: out_v[104] = 10'b0101011110;
    16'b0000001100100000: out_v[104] = 10'b1111000011;
    16'b0000010100100000: out_v[104] = 10'b0101011000;
    16'b0000001100110000: out_v[104] = 10'b1111100110;
    16'b0000011000100000: out_v[104] = 10'b0011010010;
    16'b0001000100000100: out_v[104] = 10'b1101100101;
    16'b0000000100000100: out_v[104] = 10'b0011000101;
    16'b0000011100010101: out_v[104] = 10'b1010100000;
    16'b0000001100010101: out_v[104] = 10'b1111001100;
    default: out_v[104] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001001000000100: out_v[105] = 10'b0010100100;
    16'b0000011000010100: out_v[105] = 10'b0001010111;
    16'b0001011000010000: out_v[105] = 10'b1101010010;
    16'b0000011000010000: out_v[105] = 10'b1101011010;
    16'b0001010000010001: out_v[105] = 10'b1000100111;
    16'b0000011000010001: out_v[105] = 10'b0111011101;
    16'b0001010000000000: out_v[105] = 10'b0011000101;
    16'b0001010000010000: out_v[105] = 10'b1100000110;
    16'b0001011000000000: out_v[105] = 10'b0100111101;
    16'b0001011000010101: out_v[105] = 10'b0110111101;
    16'b0000011000000101: out_v[105] = 10'b1100000111;
    16'b0000011000010101: out_v[105] = 10'b0101000101;
    16'b0001001000000000: out_v[105] = 10'b1001100011;
    16'b0001011000000001: out_v[105] = 10'b0010110111;
    16'b0000011000000000: out_v[105] = 10'b1110100001;
    16'b0001011000010100: out_v[105] = 10'b0000101111;
    16'b0001011000000101: out_v[105] = 10'b0110010010;
    16'b0001010000000001: out_v[105] = 10'b1000110100;
    16'b0000010000000000: out_v[105] = 10'b0111000101;
    16'b0001011000000100: out_v[105] = 10'b0101110100;
    16'b0001011000010001: out_v[105] = 10'b1111111000;
    16'b0000011000000100: out_v[105] = 10'b1000111100;
    16'b0000011100010101: out_v[105] = 10'b0010100111;
    16'b0001001000000101: out_v[105] = 10'b0011001100;
    16'b0001000000000000: out_v[105] = 10'b1110100010;
    16'b0001001000000001: out_v[105] = 10'b1010001001;
    16'b0001001000010101: out_v[105] = 10'b1110111001;
    16'b0000010000010000: out_v[105] = 10'b0110101101;
    16'b0000001000000000: out_v[105] = 10'b1000111011;
    16'b0000010000000001: out_v[105] = 10'b0111011100;
    16'b0000000000000001: out_v[105] = 10'b1001001111;
    16'b0000000000000000: out_v[105] = 10'b0011011010;
    16'b0000000000010000: out_v[105] = 10'b0111001101;
    16'b0000000000010001: out_v[105] = 10'b0011010111;
    16'b0001000000010000: out_v[105] = 10'b0010011110;
    16'b0000000000000101: out_v[105] = 10'b1100010101;
    16'b0001000000010101: out_v[105] = 10'b0100011011;
    16'b0001000000010001: out_v[105] = 10'b0000011110;
    16'b0000000000010101: out_v[105] = 10'b1000100011;
    16'b0000010000000101: out_v[105] = 10'b1001001011;
    16'b0000010000010001: out_v[105] = 10'b0101111100;
    16'b0000110000000001: out_v[105] = 10'b1010001010;
    16'b0001000000000001: out_v[105] = 10'b1110001100;
    16'b0000001000000100: out_v[105] = 10'b0011100100;
    16'b0000111000010000: out_v[105] = 10'b1110100100;
    16'b0000111000010101: out_v[105] = 10'b1110010100;
    16'b0000001000000101: out_v[105] = 10'b0110110000;
    16'b0000111000010100: out_v[105] = 10'b0010000111;
    16'b0001110000010000: out_v[105] = 10'b0011100110;
    16'b0000111000000101: out_v[105] = 10'b0000101101;
    16'b0000010000010101: out_v[105] = 10'b0010110010;
    16'b0001111000010101: out_v[105] = 10'b1010110110;
    16'b0000110000010000: out_v[105] = 10'b1000001011;
    16'b0001111000010100: out_v[105] = 10'b0110111111;
    16'b0001010000010101: out_v[105] = 10'b1011001010;
    16'b0000110000010001: out_v[105] = 10'b0100011011;
    16'b0000111000000100: out_v[105] = 10'b1001010110;
    16'b0000001000010101: out_v[105] = 10'b1000111111;
    16'b0001110000010001: out_v[105] = 10'b1111101010;
    16'b0001111000010000: out_v[105] = 10'b0111000000;
    16'b0000011000000001: out_v[105] = 10'b1100011110;
    16'b0001000000000101: out_v[105] = 10'b1100011001;
    16'b0000110000010101: out_v[105] = 10'b1010011011;
    16'b0001010000000101: out_v[105] = 10'b1101001001;
    16'b0000000000000100: out_v[105] = 10'b0100110011;
    16'b1001001000000101: out_v[105] = 10'b0000101110;
    16'b1001000000000101: out_v[105] = 10'b1101001101;
    16'b0000010000000100: out_v[105] = 10'b1110101010;
    16'b0001000000000100: out_v[105] = 10'b1100110110;
    16'b0001010000010100: out_v[105] = 10'b1011111111;
    16'b0000001000000001: out_v[105] = 10'b0110011011;
    16'b0001000000010100: out_v[105] = 10'b1001000011;
    16'b0001001000010100: out_v[105] = 10'b1010000011;
    16'b0001001100010100: out_v[105] = 10'b0001111111;
    16'b1001001000010100: out_v[105] = 10'b1001011100;
    16'b0001001000010000: out_v[105] = 10'b1100110111;
    16'b0001001000010001: out_v[105] = 10'b1110001011;
    16'b0000001000010000: out_v[105] = 10'b1101101010;
    16'b0000001100000100: out_v[105] = 10'b1000111010;
    16'b1000001000010101: out_v[105] = 10'b0111010111;
    16'b0000001000010001: out_v[105] = 10'b1101010000;
    16'b0000001000010100: out_v[105] = 10'b0011111010;
    16'b1001001000010101: out_v[105] = 10'b1110100011;
    16'b0000001100010100: out_v[105] = 10'b1000111011;
    16'b0001001100010000: out_v[105] = 10'b0001010011;
    16'b0001010000000100: out_v[105] = 10'b0100110001;
    16'b0000010100010100: out_v[105] = 10'b1111011110;
    16'b0001011100010101: out_v[105] = 10'b1010100010;
    16'b0001010100010100: out_v[105] = 10'b1011001111;
    16'b0000010100010000: out_v[105] = 10'b0011011001;
    16'b0000011100010100: out_v[105] = 10'b1010111110;
    16'b0001001100010101: out_v[105] = 10'b1000111010;
    16'b0001011100010100: out_v[105] = 10'b0110110010;
    16'b0001011100000100: out_v[105] = 10'b1001001001;
    16'b0000011100000101: out_v[105] = 10'b1011011011;
    16'b0000010100010101: out_v[105] = 10'b1100110011;
    16'b1001001000000100: out_v[105] = 10'b0011100111;
    16'b0000010100000101: out_v[105] = 10'b1101111000;
    16'b0001001100000100: out_v[105] = 10'b1111100000;
    16'b0000001100010101: out_v[105] = 10'b0111001111;
    16'b0001010100000100: out_v[105] = 10'b1001110110;
    16'b0000010000010100: out_v[105] = 10'b0110100110;
    16'b0001010100010101: out_v[105] = 10'b1001110011;
    16'b0000000000010100: out_v[105] = 10'b1001001100;
    16'b0001101000010100: out_v[105] = 10'b1110111110;
    16'b0000100000000100: out_v[105] = 10'b1001000001;
    16'b0000101000000100: out_v[105] = 10'b1111100001;
    16'b0001100000000100: out_v[105] = 10'b1111011101;
    16'b0001101000000100: out_v[105] = 10'b1100111011;
    16'b0001101000010000: out_v[105] = 10'b0011011000;
    16'b0001100000010100: out_v[105] = 10'b1011011011;
    16'b0000101000010100: out_v[105] = 10'b1110100111;
    16'b0001101000000000: out_v[105] = 10'b0101001111;
    16'b0000100000010100: out_v[105] = 10'b1011010000;
    16'b0001111000000000: out_v[105] = 10'b1111000010;
    16'b0001111000000100: out_v[105] = 10'b0011011111;
    16'b1001000000000001: out_v[105] = 10'b0101010101;
    16'b1001000000010001: out_v[105] = 10'b0010110001;
    16'b1001000000010000: out_v[105] = 10'b1110101000;
    16'b1000000000010001: out_v[105] = 10'b0011100011;
    16'b1001001000010001: out_v[105] = 10'b1010110100;
    16'b1000000000000001: out_v[105] = 10'b0100111010;
    16'b1001001000000001: out_v[105] = 10'b1100111110;
    16'b1001000000010101: out_v[105] = 10'b1111100101;
    16'b1001001000010000: out_v[105] = 10'b0011100001;
    16'b1001001000000000: out_v[105] = 10'b1001101011;
    default: out_v[105] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100000000000100: out_v[106] = 10'b0111010101;
    16'b1100000000000110: out_v[106] = 10'b1001111001;
    16'b1100000000000010: out_v[106] = 10'b0010111101;
    16'b1101010000010010: out_v[106] = 10'b1111010111;
    16'b1101000000000110: out_v[106] = 10'b1011101011;
    16'b0100010000000000: out_v[106] = 10'b0111011011;
    16'b1100010000000010: out_v[106] = 10'b0001110001;
    16'b0000010000000000: out_v[106] = 10'b1100010001;
    16'b1101000000010100: out_v[106] = 10'b1110001011;
    16'b1100000000000100: out_v[106] = 10'b0100111001;
    16'b0100000000000110: out_v[106] = 10'b0011001101;
    16'b1100000000010110: out_v[106] = 10'b1010100111;
    16'b1101000000000010: out_v[106] = 10'b0101110101;
    16'b1101010000010110: out_v[106] = 10'b1101100111;
    16'b0101000000000110: out_v[106] = 10'b1111001100;
    16'b1100010000000110: out_v[106] = 10'b0101011011;
    16'b1101000000010110: out_v[106] = 10'b1011011001;
    16'b0100010000010000: out_v[106] = 10'b1001011111;
    16'b1100000000000000: out_v[106] = 10'b0011100000;
    16'b1101000000010010: out_v[106] = 10'b0101101110;
    16'b1100010000000000: out_v[106] = 10'b0110110110;
    16'b1100000000010100: out_v[106] = 10'b0110010010;
    16'b0101010000010010: out_v[106] = 10'b1110111001;
    16'b1101000000000100: out_v[106] = 10'b1001110011;
    16'b0100010000000010: out_v[106] = 10'b0001010111;
    16'b1100010000010010: out_v[106] = 10'b0011011011;
    16'b0100010000010010: out_v[106] = 10'b0110110111;
    16'b0000010000000010: out_v[106] = 10'b1101101011;
    16'b0101010000010000: out_v[106] = 10'b1011011011;
    16'b0100000000000000: out_v[106] = 10'b0101110110;
    16'b1000000000000110: out_v[106] = 10'b1101010000;
    16'b0101000000000100: out_v[106] = 10'b1111100111;
    16'b1101010000010000: out_v[106] = 10'b1010011110;
    16'b1000000000000010: out_v[106] = 10'b1101010110;
    16'b0101000000010110: out_v[106] = 10'b1110100100;
    16'b1101000000010000: out_v[106] = 10'b1111011001;
    16'b0000000000000000: out_v[106] = 10'b0000110100;
    16'b0001000000000000: out_v[106] = 10'b0111011001;
    16'b0000000000010000: out_v[106] = 10'b1111100010;
    16'b0101000000000000: out_v[106] = 10'b0000101010;
    16'b0000000000000100: out_v[106] = 10'b0010101111;
    16'b0001000000010000: out_v[106] = 10'b0110100010;
    16'b0101000000010000: out_v[106] = 10'b0001101110;
    16'b0000000000011000: out_v[106] = 10'b1000001001;
    16'b0000000000000110: out_v[106] = 10'b0001101100;
    16'b0101000000010100: out_v[106] = 10'b0110000100;
    16'b0001000000000100: out_v[106] = 10'b0001011000;
    16'b0001000000010100: out_v[106] = 10'b1101001011;
    16'b1000000000000100: out_v[106] = 10'b1001100010;
    16'b0100100000011000: out_v[106] = 10'b0001111111;
    16'b0000000000010100: out_v[106] = 10'b0010111001;
    16'b0101000000011000: out_v[106] = 10'b0110111001;
    16'b0101100000011000: out_v[106] = 10'b1000100110;
    16'b0100000000010000: out_v[106] = 10'b0111100010;
    16'b1001000000000100: out_v[106] = 10'b0010010101;
    16'b0101000000001000: out_v[106] = 10'b0111011111;
    16'b0100000000011000: out_v[106] = 10'b1100010000;
    16'b0001000000000110: out_v[106] = 10'b1110010110;
    16'b0101000000011100: out_v[106] = 10'b1001010111;
    16'b0000000000010110: out_v[106] = 10'b1100110110;
    16'b0001000000010110: out_v[106] = 10'b1011010101;
    16'b0000000000011100: out_v[106] = 10'b0110001111;
    16'b0101000000011110: out_v[106] = 10'b1111010010;
    16'b0000100000011000: out_v[106] = 10'b1001010101;
    16'b0100000000010100: out_v[106] = 10'b0100001110;
    16'b1001000000010100: out_v[106] = 10'b0111001111;
    16'b0001000000011100: out_v[106] = 10'b1011111010;
    16'b0101000000000010: out_v[106] = 10'b0010111000;
    16'b0100000000010010: out_v[106] = 10'b1110111000;
    16'b0101000000001010: out_v[106] = 10'b0100011001;
    16'b0100000000011110: out_v[106] = 10'b1111100100;
    16'b1100000000011010: out_v[106] = 10'b0011010111;
    16'b0000100000011010: out_v[106] = 10'b1101000010;
    16'b0100000000011010: out_v[106] = 10'b1010011011;
    16'b0100100000011010: out_v[106] = 10'b1101100100;
    16'b0100000000000010: out_v[106] = 10'b1111001010;
    16'b0100000010000000: out_v[106] = 10'b1010000001;
    16'b0101000000011010: out_v[106] = 10'b0011101010;
    16'b0000000000011010: out_v[106] = 10'b1100001010;
    16'b0101000000010010: out_v[106] = 10'b0000110011;
    16'b0000000000010010: out_v[106] = 10'b0101100001;
    16'b0100000010010000: out_v[106] = 10'b1111111010;
    16'b1000000000001110: out_v[106] = 10'b0001011011;
    16'b0000010000000110: out_v[106] = 10'b1100110011;
    16'b1000000000000000: out_v[106] = 10'b0101011110;
    16'b1000000000010000: out_v[106] = 10'b0011001101;
    16'b1000000000010100: out_v[106] = 10'b1110110100;
    16'b1000010000000100: out_v[106] = 10'b0110111100;
    16'b1000000000010110: out_v[106] = 10'b1100100111;
    16'b1000010000000110: out_v[106] = 10'b1110010011;
    16'b1000110000001110: out_v[106] = 10'b1000011110;
    16'b1000000000001100: out_v[106] = 10'b0011011111;
    16'b1000010000000000: out_v[106] = 10'b0110101101;
    16'b1000010000010110: out_v[106] = 10'b0100110000;
    16'b1100010000000100: out_v[106] = 10'b0101011111;
    16'b0000010000000100: out_v[106] = 10'b1000000001;
    16'b1100000000010010: out_v[106] = 10'b0011101110;
    16'b0100000100000000: out_v[106] = 10'b0100100001;
    16'b0100000000010110: out_v[106] = 10'b1110100011;
    16'b1100000000010000: out_v[106] = 10'b0111010110;
    16'b1001000000010110: out_v[106] = 10'b0111011000;
    16'b0001000000000010: out_v[106] = 10'b1101101000;
    16'b1001000000000110: out_v[106] = 10'b1100010111;
    16'b0100100000000000: out_v[106] = 10'b1100011111;
    16'b0000100000001010: out_v[106] = 10'b0010001100;
    16'b0000100000000000: out_v[106] = 10'b0100111011;
    16'b0000100000001000: out_v[106] = 10'b1110000110;
    16'b0000000000001000: out_v[106] = 10'b1010010010;
    16'b0100000000001000: out_v[106] = 10'b0011010011;
    16'b0000100000000010: out_v[106] = 10'b1001010111;
    16'b0000100001000000: out_v[106] = 10'b1001011100;
    16'b0100100000001000: out_v[106] = 10'b1011010011;
    16'b1000000001000100: out_v[106] = 10'b1101001011;
    default: out_v[106] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100000000000000: out_v[107] = 10'b1111000001;
    16'b0100000000000010: out_v[107] = 10'b1100011000;
    16'b0100010000000000: out_v[107] = 10'b1111000011;
    16'b1000000000000010: out_v[107] = 10'b1010101111;
    16'b0000000000000000: out_v[107] = 10'b0110100010;
    16'b0100000010000000: out_v[107] = 10'b1001011110;
    16'b0000000000000010: out_v[107] = 10'b1000011001;
    16'b1100000000000000: out_v[107] = 10'b1010010000;
    16'b0000010000000000: out_v[107] = 10'b0100100100;
    16'b0100010010000000: out_v[107] = 10'b1101011001;
    16'b1100000000000010: out_v[107] = 10'b0001010101;
    16'b1000000000000000: out_v[107] = 10'b1110110010;
    16'b1000000010000000: out_v[107] = 10'b1001001010;
    16'b1000010010000000: out_v[107] = 10'b0101110111;
    16'b0000000010000000: out_v[107] = 10'b0011110101;
    16'b0000010010000000: out_v[107] = 10'b0010100010;
    16'b1100010010000000: out_v[107] = 10'b0101010100;
    16'b1100010000000010: out_v[107] = 10'b1011011100;
    16'b1100000010000010: out_v[107] = 10'b0100010001;
    16'b1100000010000000: out_v[107] = 10'b0001010110;
    16'b1100010000000000: out_v[107] = 10'b1001001110;
    16'b1000010000000000: out_v[107] = 10'b1001000110;
    16'b0000000010000010: out_v[107] = 10'b1100100010;
    16'b0000000000100000: out_v[107] = 10'b0110011100;
    16'b0000010000100000: out_v[107] = 10'b1000001010;
    16'b0000001000000000: out_v[107] = 10'b1110101110;
    16'b0100001000000000: out_v[107] = 10'b1110100000;
    16'b1000001000000000: out_v[107] = 10'b0010010111;
    16'b1100001000000000: out_v[107] = 10'b1011110110;
    16'b1000000000010000: out_v[107] = 10'b1111100111;
    16'b0000000000010000: out_v[107] = 10'b1000011111;
    16'b1000000000100000: out_v[107] = 10'b0010011111;
    16'b1000100000000000: out_v[107] = 10'b1010011001;
    default: out_v[107] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000001000100000: out_v[108] = 10'b1100111001;
    16'b1000001000100110: out_v[108] = 10'b0111000011;
    16'b1000011000000110: out_v[108] = 10'b1101000101;
    16'b0000000000000110: out_v[108] = 10'b0101011010;
    16'b0000001000000110: out_v[108] = 10'b1110001011;
    16'b0000011000000110: out_v[108] = 10'b1000011011;
    16'b1000000000000010: out_v[108] = 10'b1001010110;
    16'b0000001000000010: out_v[108] = 10'b0001010111;
    16'b0000010000000100: out_v[108] = 10'b1001000011;
    16'b0000001000100100: out_v[108] = 10'b0110110011;
    16'b1000001000000010: out_v[108] = 10'b1000001111;
    16'b0000001000100110: out_v[108] = 10'b0100110111;
    16'b1000011000100110: out_v[108] = 10'b0100011100;
    16'b1000001000000110: out_v[108] = 10'b0100011111;
    16'b0000001000000100: out_v[108] = 10'b1010010111;
    16'b1000000000000110: out_v[108] = 10'b0010100010;
    16'b0000000000100110: out_v[108] = 10'b1101010110;
    16'b0000011000100110: out_v[108] = 10'b1110000111;
    16'b0000011000000100: out_v[108] = 10'b0011110101;
    16'b1000011000000000: out_v[108] = 10'b1100010111;
    16'b1000101000100110: out_v[108] = 10'b1011001010;
    16'b1000101000100100: out_v[108] = 10'b0011001011;
    16'b0000000000000100: out_v[108] = 10'b1101100001;
    16'b1000011000000010: out_v[108] = 10'b0100001101;
    16'b0000010000000110: out_v[108] = 10'b0111110000;
    16'b1000010000000010: out_v[108] = 10'b0111110000;
    16'b1000001000100100: out_v[108] = 10'b1010001011;
    16'b1000010000000110: out_v[108] = 10'b0100111100;
    16'b0000011000000010: out_v[108] = 10'b1100001011;
    16'b1000001000100010: out_v[108] = 10'b1000001110;
    16'b1000101000000010: out_v[108] = 10'b1001110000;
    16'b0000000000100100: out_v[108] = 10'b1000110000;
    16'b1000011000000100: out_v[108] = 10'b1001010111;
    16'b0000001000100010: out_v[108] = 10'b1101010000;
    16'b0000101000000000: out_v[108] = 10'b0101000101;
    16'b0000001000000000: out_v[108] = 10'b1110001010;
    16'b0000000000000000: out_v[108] = 10'b1110100011;
    16'b1000101000000100: out_v[108] = 10'b1100111001;
    16'b1000001000000100: out_v[108] = 10'b0111010100;
    16'b0000101000000100: out_v[108] = 10'b1110110010;
    16'b0000000000100000: out_v[108] = 10'b1001110000;
    16'b0000011000000000: out_v[108] = 10'b1011000101;
    16'b1000000000000100: out_v[108] = 10'b0100010111;
    16'b0000010000000000: out_v[108] = 10'b1000100110;
    16'b1000010000000100: out_v[108] = 10'b0010110111;
    16'b0000000000000010: out_v[108] = 10'b0111110100;
    16'b0000011000100100: out_v[108] = 10'b0110010111;
    16'b1000110000000100: out_v[108] = 10'b0011100101;
    16'b1000100000000100: out_v[108] = 10'b0011000101;
    16'b1000010000000000: out_v[108] = 10'b0011101011;
    16'b0000010000000010: out_v[108] = 10'b1101100010;
    16'b1000000000000000: out_v[108] = 10'b0001101001;
    16'b1000001000000000: out_v[108] = 10'b0011111011;
    16'b1000111000000100: out_v[108] = 10'b1011100101;
    16'b1000001000100000: out_v[108] = 10'b1110110000;
    16'b0000001010000000: out_v[108] = 10'b0011101001;
    16'b1000010000100010: out_v[108] = 10'b0000111100;
    16'b0000011000100010: out_v[108] = 10'b0001101001;
    16'b0000011010100010: out_v[108] = 10'b1000001111;
    16'b0000000000100010: out_v[108] = 10'b0000100010;
    16'b0000011000100000: out_v[108] = 10'b1010011000;
    16'b1000011000100010: out_v[108] = 10'b1001000100;
    16'b0000010000100010: out_v[108] = 10'b1010111001;
    16'b1000000000100010: out_v[108] = 10'b1011100100;
    16'b0000001010100000: out_v[108] = 10'b1100100010;
    16'b0000011000110010: out_v[108] = 10'b1001101100;
    16'b1000000000100000: out_v[108] = 10'b1001101110;
    16'b0000000010100000: out_v[108] = 10'b0000010111;
    16'b0100001000100000: out_v[108] = 10'b0100011110;
    16'b0000000010000000: out_v[108] = 10'b0110111011;
    16'b0000100000000100: out_v[108] = 10'b1110010100;
    16'b0000100000000000: out_v[108] = 10'b0110100010;
    16'b0000100000000110: out_v[108] = 10'b0101011110;
    16'b0000100000100000: out_v[108] = 10'b1111011101;
    16'b0100001000000000: out_v[108] = 10'b1011000111;
    16'b0000100000100100: out_v[108] = 10'b1101001010;
    16'b0001001000100100: out_v[108] = 10'b0111001110;
    16'b0001001000000000: out_v[108] = 10'b1110110111;
    16'b0000010000100110: out_v[108] = 10'b1011010000;
    16'b0000010000100000: out_v[108] = 10'b0100100011;
    16'b1000110000100010: out_v[108] = 10'b1100100100;
    16'b0001001000100000: out_v[108] = 10'b1010100101;
    16'b1000101000100000: out_v[108] = 10'b0010101110;
    16'b0000101000100100: out_v[108] = 10'b0011000010;
    16'b0000111000100110: out_v[108] = 10'b1011000010;
    16'b0000101000100110: out_v[108] = 10'b1101000111;
    16'b0000110000000110: out_v[108] = 10'b1101011010;
    16'b0000001010000010: out_v[108] = 10'b1010000010;
    16'b0100001000000010: out_v[108] = 10'b0111000011;
    16'b0100011000000010: out_v[108] = 10'b0010101111;
    16'b0100001100000000: out_v[108] = 10'b1001111110;
    16'b0000001110000000: out_v[108] = 10'b0110110110;
    16'b0100000000000000: out_v[108] = 10'b1111001010;
    16'b0000001100000000: out_v[108] = 10'b1001111100;
    16'b1000000000100100: out_v[108] = 10'b1011001011;
    16'b0000001010000100: out_v[108] = 10'b0000011010;
    16'b0100001000000100: out_v[108] = 10'b1101101010;
    16'b0100011000000110: out_v[108] = 10'b1000110110;
    16'b0100011000000000: out_v[108] = 10'b0111111000;
    16'b0100000000100000: out_v[108] = 10'b0001011101;
    default: out_v[108] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000000000010: out_v[109] = 10'b1111000011;
    16'b0001000000000001: out_v[109] = 10'b1000001001;
    16'b0001000000000010: out_v[109] = 10'b0101100001;
    16'b0000000000000110: out_v[109] = 10'b1110010010;
    16'b0000000000000000: out_v[109] = 10'b1110000110;
    16'b0001000001001101: out_v[109] = 10'b0000111111;
    16'b0001000000000000: out_v[109] = 10'b1011100000;
    16'b0001000000000011: out_v[109] = 10'b0111010000;
    16'b0001000001000001: out_v[109] = 10'b1011011111;
    16'b0001000000000110: out_v[109] = 10'b1001100011;
    16'b0001000000000101: out_v[109] = 10'b0000101101;
    16'b0000000000000001: out_v[109] = 10'b0001101011;
    16'b0001000001001001: out_v[109] = 10'b1000001001;
    16'b0001000001000111: out_v[109] = 10'b0100111111;
    16'b0001000000000111: out_v[109] = 10'b0111100000;
    16'b0001000001000000: out_v[109] = 10'b0010000111;
    16'b0001000000000100: out_v[109] = 10'b1101110110;
    16'b0001000001000101: out_v[109] = 10'b1011001111;
    16'b0000000000000100: out_v[109] = 10'b1010101110;
    16'b0000000000000111: out_v[109] = 10'b0101000010;
    16'b0001000001000011: out_v[109] = 10'b1110010111;
    16'b0011000000000001: out_v[109] = 10'b0111010101;
    16'b0000000000000011: out_v[109] = 10'b1001000110;
    16'b0001000001001111: out_v[109] = 10'b1101110101;
    16'b0000000100000000: out_v[109] = 10'b1000111110;
    16'b0000000000000101: out_v[109] = 10'b1100001110;
    16'b0000000100000110: out_v[109] = 10'b1110110111;
    16'b0000000100000010: out_v[109] = 10'b0000001111;
    16'b0000000100000101: out_v[109] = 10'b0010011101;
    16'b0000000100000100: out_v[109] = 10'b1011111100;
    16'b0001000001000110: out_v[109] = 10'b1111010000;
    16'b0001000001000100: out_v[109] = 10'b1110010011;
    16'b0011000001000101: out_v[109] = 10'b1010001110;
    16'b0010000000000001: out_v[109] = 10'b0111011011;
    16'b0000000100000001: out_v[109] = 10'b0100100100;
    16'b0010000000000101: out_v[109] = 10'b0011110000;
    16'b0011000000000101: out_v[109] = 10'b0001110101;
    16'b0010000100000101: out_v[109] = 10'b1001011111;
    16'b0011000000000100: out_v[109] = 10'b1100000010;
    16'b0001000100000101: out_v[109] = 10'b0000001111;
    16'b0010000000000100: out_v[109] = 10'b1100001010;
    16'b0001000001001100: out_v[109] = 10'b0101010100;
    16'b0001000000001100: out_v[109] = 10'b0111001100;
    16'b0001000100000110: out_v[109] = 10'b1110110111;
    16'b0001000001001110: out_v[109] = 10'b0000111010;
    16'b0001000000001110: out_v[109] = 10'b0001011111;
    16'b0000000001001100: out_v[109] = 10'b1100101010;
    16'b0000000001001001: out_v[109] = 10'b0110110110;
    16'b0011000001001101: out_v[109] = 10'b0100110101;
    16'b0000000001001101: out_v[109] = 10'b0110110010;
    16'b0001000001001010: out_v[109] = 10'b1000101000;
    16'b0000000001000001: out_v[109] = 10'b1111110110;
    16'b0001000001001000: out_v[109] = 10'b1010101101;
    16'b0000000001000100: out_v[109] = 10'b1000100111;
    16'b0000000001000101: out_v[109] = 10'b0111000110;
    16'b0000000001000000: out_v[109] = 10'b0001101001;
    16'b0000000001001000: out_v[109] = 10'b1010111100;
    16'b0100000000000110: out_v[109] = 10'b1010101110;
    16'b0001000100000100: out_v[109] = 10'b1010101011;
    16'b0011000001001011: out_v[109] = 10'b0000010110;
    16'b0001000001001011: out_v[109] = 10'b1011000111;
    16'b0001000001000010: out_v[109] = 10'b0100001100;
    default: out_v[109] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010000001001010: out_v[110] = 10'b1100001111;
    16'b0011000001001000: out_v[110] = 10'b1100011010;
    16'b0011000001000000: out_v[110] = 10'b0010101101;
    16'b0000000001001010: out_v[110] = 10'b1101010011;
    16'b0000001001001010: out_v[110] = 10'b0010110010;
    16'b0010001001001000: out_v[110] = 10'b0110000101;
    16'b0010000000001000: out_v[110] = 10'b0100100011;
    16'b0010000001000000: out_v[110] = 10'b1101000011;
    16'b0010100001000000: out_v[110] = 10'b1111000011;
    16'b0000001000001010: out_v[110] = 10'b0011011011;
    16'b0011000001001010: out_v[110] = 10'b0100110001;
    16'b0000000000000010: out_v[110] = 10'b0010100110;
    16'b0000100100000000: out_v[110] = 10'b0111100101;
    16'b0010000001000010: out_v[110] = 10'b1101000011;
    16'b0011001001001000: out_v[110] = 10'b0001110011;
    16'b0001001001001000: out_v[110] = 10'b1011001011;
    16'b0010100001001000: out_v[110] = 10'b0111110011;
    16'b0000000001000000: out_v[110] = 10'b0010010000;
    16'b0000000000001010: out_v[110] = 10'b0011011010;
    16'b0010100101000000: out_v[110] = 10'b1001000001;
    16'b0000100101000000: out_v[110] = 10'b1000101011;
    16'b0010100101001010: out_v[110] = 10'b1000010101;
    16'b0010001001001010: out_v[110] = 10'b1110101011;
    16'b0000000001000010: out_v[110] = 10'b0010001111;
    16'b0000100101000010: out_v[110] = 10'b0101011011;
    16'b0011000000001000: out_v[110] = 10'b0110110111;
    16'b0010100101001000: out_v[110] = 10'b1010011011;
    16'b0010100101000010: out_v[110] = 10'b1010011011;
    16'b0000000000001000: out_v[110] = 10'b1100100001;
    16'b0011100001000000: out_v[110] = 10'b1111011111;
    16'b0010000001001000: out_v[110] = 10'b1011111110;
    16'b0010100001001010: out_v[110] = 10'b1010001011;
    16'b0001001001001010: out_v[110] = 10'b1110011111;
    16'b0000000001001000: out_v[110] = 10'b0101010011;
    16'b0001000001001000: out_v[110] = 10'b0100110010;
    16'b0000001001000000: out_v[110] = 10'b0010001011;
    16'b0011100101000000: out_v[110] = 10'b1110000001;
    16'b0000001000000010: out_v[110] = 10'b0110100010;
    16'b0011001001001010: out_v[110] = 10'b0010001001;
    16'b0000001001001000: out_v[110] = 10'b1001110010;
    16'b0000001001000010: out_v[110] = 10'b1110010000;
    16'b0011100101001000: out_v[110] = 10'b0101011011;
    16'b0000001000001000: out_v[110] = 10'b0000101001;
    16'b0000000000000000: out_v[110] = 10'b0111100011;
    16'b0011001001000000: out_v[110] = 10'b1001110001;
    16'b0011100001001000: out_v[110] = 10'b1111010111;
    16'b0010100001000010: out_v[110] = 10'b0111111111;
    16'b0000100000000000: out_v[110] = 10'b1101000111;
    16'b0000100100000010: out_v[110] = 10'b0110101101;
    16'b0001000001000000: out_v[110] = 10'b1100011010;
    16'b0000000100001000: out_v[110] = 10'b0010110010;
    16'b0000000100000000: out_v[110] = 10'b1001100100;
    16'b0000100001000010: out_v[110] = 10'b0010101100;
    16'b0000001000000000: out_v[110] = 10'b0010100100;
    16'b0001100000000000: out_v[110] = 10'b0101011011;
    16'b0000101000000010: out_v[110] = 10'b1001010011;
    16'b0000100001000000: out_v[110] = 10'b1001011010;
    16'b0000000101000000: out_v[110] = 10'b0101000110;
    16'b0001100001000000: out_v[110] = 10'b1101000111;
    16'b0000100000000010: out_v[110] = 10'b0011011011;
    16'b0000101001000000: out_v[110] = 10'b1111000100;
    16'b0001100001000010: out_v[110] = 10'b1101101001;
    16'b0011101001000010: out_v[110] = 10'b0110111100;
    16'b0001101001000010: out_v[110] = 10'b1110110011;
    16'b0001001001000000: out_v[110] = 10'b0101011100;
    16'b0000101001000010: out_v[110] = 10'b0011110011;
    16'b0001000001000010: out_v[110] = 10'b1001001110;
    16'b0001101000000010: out_v[110] = 10'b0001000101;
    16'b0000100000001000: out_v[110] = 10'b1010111111;
    16'b0000101000000000: out_v[110] = 10'b1101001110;
    16'b0001001001000010: out_v[110] = 10'b1011110110;
    16'b0001101001000000: out_v[110] = 10'b0100000101;
    16'b0000100000001010: out_v[110] = 10'b0111110100;
    16'b0001000101000000: out_v[110] = 10'b1000110111;
    16'b0011001001000010: out_v[110] = 10'b1011110110;
    16'b0001001000001000: out_v[110] = 10'b0011101100;
    16'b0001001000000000: out_v[110] = 10'b0100011101;
    16'b1000101100001000: out_v[110] = 10'b1001001011;
    16'b0000001100001000: out_v[110] = 10'b0011111011;
    16'b0000001100000000: out_v[110] = 10'b1000010100;
    16'b0000100100001000: out_v[110] = 10'b0000101100;
    16'b0000101100001000: out_v[110] = 10'b1010011010;
    16'b1000100100001000: out_v[110] = 10'b0011001000;
    16'b0000101100000000: out_v[110] = 10'b0010111011;
    16'b0000101000001000: out_v[110] = 10'b0011011111;
    16'b0001000000001000: out_v[110] = 10'b0111110000;
    16'b0001100001001000: out_v[110] = 10'b1011111000;
    16'b0001000000000000: out_v[110] = 10'b1110000011;
    16'b0000001100000010: out_v[110] = 10'b0001111011;
    16'b0000001101000010: out_v[110] = 10'b0010010011;
    16'b0000000100000010: out_v[110] = 10'b0011011011;
    16'b0000001101000000: out_v[110] = 10'b0110010111;
    16'b0000001101001010: out_v[110] = 10'b1001011011;
    16'b0000001100001010: out_v[110] = 10'b0111011001;
    16'b0010001000001010: out_v[110] = 10'b0011011010;
    16'b0010001001000010: out_v[110] = 10'b1000111010;
    16'b0000001101001000: out_v[110] = 10'b0001110110;
    16'b0000000101001000: out_v[110] = 10'b1100001110;
    16'b0000100101001000: out_v[110] = 10'b0000100110;
    16'b0000101000001010: out_v[110] = 10'b1011001110;
    16'b0010100000000000: out_v[110] = 10'b0011111000;
    16'b0010100000000010: out_v[110] = 10'b1010111111;
    16'b0010000000000010: out_v[110] = 10'b0101001100;
    16'b0010000000001010: out_v[110] = 10'b1011011011;
    16'b0010001000000010: out_v[110] = 10'b0101111110;
    16'b0010000000000000: out_v[110] = 10'b0011111000;
    16'b0010001001000000: out_v[110] = 10'b1011100010;
    16'b0010001000001000: out_v[110] = 10'b0110110111;
    16'b0000000101001010: out_v[110] = 10'b1110000000;
    16'b0000101101001000: out_v[110] = 10'b0111010101;
    16'b0001000001001010: out_v[110] = 10'b0100000111;
    16'b0000101101000000: out_v[110] = 10'b0111111011;
    16'b0000100100001010: out_v[110] = 10'b1100000110;
    16'b0000101101001010: out_v[110] = 10'b0101110010;
    default: out_v[110] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0101100010000100: out_v[111] = 10'b1110001011;
    16'b0101000010010100: out_v[111] = 10'b0101000011;
    16'b0000100010110100: out_v[111] = 10'b0110110011;
    16'b0101000010000100: out_v[111] = 10'b0111011000;
    16'b0001000010110000: out_v[111] = 10'b0001010011;
    16'b0000100010110000: out_v[111] = 10'b1111110001;
    16'b0111100010010100: out_v[111] = 10'b0100100111;
    16'b0001100010110000: out_v[111] = 10'b1000110011;
    16'b0001100010010100: out_v[111] = 10'b1111101011;
    16'b0000100010000100: out_v[111] = 10'b1001000111;
    16'b0001000000110000: out_v[111] = 10'b1100010011;
    16'b0001100010000100: out_v[111] = 10'b1100110000;
    16'b0001100010110100: out_v[111] = 10'b1010001111;
    16'b0000100010010100: out_v[111] = 10'b0001111100;
    16'b1000100110110100: out_v[111] = 10'b1010011111;
    16'b1000100110110000: out_v[111] = 10'b0001000001;
    16'b0000000010110000: out_v[111] = 10'b1111011010;
    16'b1000000100100100: out_v[111] = 10'b1000001011;
    16'b0001000010010100: out_v[111] = 10'b0001100111;
    16'b0000100110010100: out_v[111] = 10'b0111010111;
    16'b0001100010010000: out_v[111] = 10'b1000001100;
    16'b0101100010010100: out_v[111] = 10'b1000001011;
    16'b1000100110100100: out_v[111] = 10'b1111101011;
    16'b1000000110110000: out_v[111] = 10'b1110001110;
    16'b0001000010110100: out_v[111] = 10'b1001101000;
    16'b1000100110000100: out_v[111] = 10'b1011011011;
    16'b0111100010000100: out_v[111] = 10'b0111000011;
    16'b0001000010010000: out_v[111] = 10'b1001100111;
    16'b0000100010010000: out_v[111] = 10'b1101110110;
    16'b0101100010000000: out_v[111] = 10'b1001001011;
    16'b0100100010000100: out_v[111] = 10'b1101100110;
    16'b0111000010010100: out_v[111] = 10'b0011010100;
    16'b1000000110110100: out_v[111] = 10'b1110010011;
    16'b1000100110010100: out_v[111] = 10'b0001011110;
    16'b1001100110110100: out_v[111] = 10'b1011101110;
    16'b0101100010110100: out_v[111] = 10'b0011011011;
    16'b0110000010010000: out_v[111] = 10'b1010111000;
    16'b0010000010000000: out_v[111] = 10'b1101010011;
    16'b0010000000000000: out_v[111] = 10'b1100001110;
    16'b0010100000000000: out_v[111] = 10'b1001000011;
    16'b0010100010000000: out_v[111] = 10'b0000011011;
    16'b0000000000000000: out_v[111] = 10'b0100000111;
    16'b0010000000010000: out_v[111] = 10'b0100101011;
    16'b0110000010000000: out_v[111] = 10'b0011010011;
    16'b0011000000000000: out_v[111] = 10'b1101011001;
    16'b0000100000000000: out_v[111] = 10'b0100100111;
    16'b0010000010010000: out_v[111] = 10'b0110011000;
    16'b0110000000010100: out_v[111] = 10'b1101001011;
    16'b0110000000010000: out_v[111] = 10'b1010110101;
    16'b0110100010000000: out_v[111] = 10'b0010001010;
    16'b0000000010000000: out_v[111] = 10'b0111001010;
    16'b0011100000000000: out_v[111] = 10'b0110100011;
    16'b0110100010010100: out_v[111] = 10'b0110100110;
    16'b0100100010010100: out_v[111] = 10'b1100101010;
    16'b0010100010010000: out_v[111] = 10'b0001011101;
    16'b0110000000000000: out_v[111] = 10'b0111001101;
    16'b0110100010000100: out_v[111] = 10'b0111101101;
    16'b1010000100000000: out_v[111] = 10'b0000111101;
    16'b0000100110000000: out_v[111] = 10'b1011110110;
    16'b0110000010010100: out_v[111] = 10'b0101010110;
    16'b0110000010000100: out_v[111] = 10'b0101011010;
    16'b1000100110010000: out_v[111] = 10'b1000011110;
    16'b0110100110010100: out_v[111] = 10'b0010000101;
    16'b0100000010010100: out_v[111] = 10'b1000000101;
    16'b0110100010010000: out_v[111] = 10'b0000111010;
    16'b1110100110010100: out_v[111] = 10'b0100011110;
    16'b1000100110000000: out_v[111] = 10'b0010111100;
    16'b0110000000000100: out_v[111] = 10'b0101000110;
    16'b0100100000010100: out_v[111] = 10'b0010001100;
    16'b0000100010000000: out_v[111] = 10'b1110110010;
    16'b1100100110010100: out_v[111] = 10'b1111101100;
    16'b0000100110010000: out_v[111] = 10'b1010001111;
    16'b1110100110000100: out_v[111] = 10'b0001111110;
    16'b0110100000010100: out_v[111] = 10'b1110101101;
    16'b0100000000000100: out_v[111] = 10'b1000011000;
    16'b0110100110010000: out_v[111] = 10'b1011001001;
    16'b0100100110010100: out_v[111] = 10'b1110100011;
    16'b1110000100000000: out_v[111] = 10'b1010110111;
    16'b0100100010010000: out_v[111] = 10'b1000001111;
    16'b0110100110000100: out_v[111] = 10'b1100111110;
    16'b1110000100000100: out_v[111] = 10'b0011101010;
    16'b1010100110010000: out_v[111] = 10'b0110011010;
    16'b0100100010000000: out_v[111] = 10'b1101001000;
    16'b1110100110010000: out_v[111] = 10'b1011101011;
    16'b1010100110000000: out_v[111] = 10'b1011001011;
    16'b1000000100000000: out_v[111] = 10'b0100010101;
    16'b0110100110000000: out_v[111] = 10'b0001111110;
    16'b0011100010000000: out_v[111] = 10'b1110100000;
    16'b0010100110010000: out_v[111] = 10'b0111010011;
    16'b0001100010000000: out_v[111] = 10'b1000001110;
    16'b0010000100000000: out_v[111] = 10'b1001001100;
    16'b1011000100000000: out_v[111] = 10'b1110010011;
    16'b0010100110000000: out_v[111] = 10'b1010111100;
    16'b0011000100000000: out_v[111] = 10'b1100001011;
    16'b0011100010010000: out_v[111] = 10'b1111000010;
    16'b1110100110000000: out_v[111] = 10'b0011111001;
    16'b0001000000000000: out_v[111] = 10'b0111001000;
    16'b0011100110010000: out_v[111] = 10'b0000011111;
    16'b0010100010010100: out_v[111] = 10'b0010001011;
    16'b0001100000010000: out_v[111] = 10'b1101001100;
    16'b0001100000000000: out_v[111] = 10'b1000101010;
    16'b0111100010010000: out_v[111] = 10'b0010111110;
    16'b0100000010000000: out_v[111] = 10'b1000110001;
    16'b0100000000100100: out_v[111] = 10'b1000011011;
    16'b0110000110000000: out_v[111] = 10'b0110101001;
    16'b0111100000000000: out_v[111] = 10'b0011001101;
    16'b0111000000000000: out_v[111] = 10'b1001100010;
    16'b0111000000000100: out_v[111] = 10'b1010111111;
    16'b1110000100100000: out_v[111] = 10'b1001101111;
    16'b0111000010000000: out_v[111] = 10'b1000100100;
    16'b0101000000000100: out_v[111] = 10'b0010111001;
    16'b0011000000000001: out_v[111] = 10'b1000010111;
    16'b0101000000000000: out_v[111] = 10'b1001010010;
    16'b0111000010000100: out_v[111] = 10'b1011001100;
    16'b0111000000100000: out_v[111] = 10'b0011101111;
    16'b0100000100000000: out_v[111] = 10'b1011010011;
    16'b0101000010000000: out_v[111] = 10'b1100100000;
    16'b0111000000100100: out_v[111] = 10'b0110110111;
    16'b0100000010000100: out_v[111] = 10'b1101010101;
    16'b0011000010000000: out_v[111] = 10'b0100110001;
    16'b0101100000000000: out_v[111] = 10'b0000111011;
    16'b0110000000100000: out_v[111] = 10'b1111100111;
    16'b0101000000100100: out_v[111] = 10'b1100111011;
    16'b1100000100000000: out_v[111] = 10'b0001100011;
    16'b0110000000100100: out_v[111] = 10'b1001010011;
    16'b1110000110000100: out_v[111] = 10'b0010111001;
    16'b1110000100100100: out_v[111] = 10'b1101010111;
    16'b1100000100100100: out_v[111] = 10'b1000111110;
    16'b0110000100000000: out_v[111] = 10'b0111011011;
    16'b0010000000100000: out_v[111] = 10'b0111001011;
    16'b1110000110000000: out_v[111] = 10'b0000111110;
    16'b0100000000000000: out_v[111] = 10'b1100100111;
    16'b1110000110100100: out_v[111] = 10'b1000111101;
    16'b1100000110000100: out_v[111] = 10'b0010000111;
    16'b0101100000000100: out_v[111] = 10'b0110011100;
    16'b0011000000100000: out_v[111] = 10'b1110101111;
    16'b0011000010010000: out_v[111] = 10'b1110100010;
    16'b0111100010000000: out_v[111] = 10'b0011100110;
    16'b0011000000010000: out_v[111] = 10'b1001111000;
    16'b1001100110010000: out_v[111] = 10'b1111110110;
    16'b0111000010010000: out_v[111] = 10'b0010100110;
    16'b0111000000010100: out_v[111] = 10'b0111111010;
    16'b0111000000010000: out_v[111] = 10'b0110101100;
    16'b0010000000000100: out_v[111] = 10'b0001111000;
    16'b0011000000000100: out_v[111] = 10'b0100101010;
    16'b0001000010000000: out_v[111] = 10'b0011001110;
    16'b0001000000010000: out_v[111] = 10'b1011100000;
    16'b0101000000010000: out_v[111] = 10'b1101111000;
    16'b0011000010000001: out_v[111] = 10'b1001000111;
    16'b0111100000000100: out_v[111] = 10'b0011110000;
    16'b1100000100001100: out_v[111] = 10'b1110111111;
    16'b0100100000000000: out_v[111] = 10'b1011000001;
    16'b0001100000000100: out_v[111] = 10'b1001010100;
    16'b0110100000000000: out_v[111] = 10'b1100010101;
    16'b1110000100001100: out_v[111] = 10'b1100011111;
    16'b0000000000000100: out_v[111] = 10'b1101011010;
    16'b1100000100000100: out_v[111] = 10'b0111011011;
    16'b0110100000000100: out_v[111] = 10'b1100111001;
    16'b0000100000000100: out_v[111] = 10'b1111011101;
    16'b0000000110000000: out_v[111] = 10'b0011100000;
    16'b0001000000100000: out_v[111] = 10'b0110100100;
    16'b1001000100000001: out_v[111] = 10'b0111010001;
    16'b0001000000000001: out_v[111] = 10'b0110001000;
    16'b1001000100000000: out_v[111] = 10'b0110000110;
    16'b1000000000000000: out_v[111] = 10'b0100110001;
    16'b0000000000000001: out_v[111] = 10'b0010110010;
    16'b1001000000000000: out_v[111] = 10'b0000110111;
    16'b1000000100000001: out_v[111] = 10'b1100001101;
    16'b1000000100100000: out_v[111] = 10'b0111001111;
    16'b0000000100000000: out_v[111] = 10'b0100010101;
    16'b0001000010000001: out_v[111] = 10'b0010111000;
    16'b1000000110000000: out_v[111] = 10'b0011111011;
    16'b1001000100100000: out_v[111] = 10'b0011010011;
    16'b0000000010000001: out_v[111] = 10'b0111011010;
    16'b0000000100000001: out_v[111] = 10'b1101110101;
    16'b0000000110000001: out_v[111] = 10'b1101010111;
    16'b1000000110000001: out_v[111] = 10'b0001110011;
    16'b1001000000000001: out_v[111] = 10'b1111010111;
    16'b0001000000100001: out_v[111] = 10'b0111011110;
    16'b1000000000000001: out_v[111] = 10'b1110110000;
    16'b0001000100000000: out_v[111] = 10'b0010101000;
    16'b0011100110000000: out_v[111] = 10'b1101110001;
    16'b1011000110000000: out_v[111] = 10'b0101010011;
    16'b0111100110010100: out_v[111] = 10'b0111000011;
    16'b1011100110000000: out_v[111] = 10'b0101010101;
    16'b1010000110000000: out_v[111] = 10'b1111000011;
    16'b1111100110000000: out_v[111] = 10'b0010110111;
    16'b0111100110000000: out_v[111] = 10'b1101100111;
    16'b0111000010000001: out_v[111] = 10'b1001010111;
    16'b0110000010000001: out_v[111] = 10'b0101100011;
    16'b0111000000000001: out_v[111] = 10'b1001100110;
    16'b0100000010100100: out_v[111] = 10'b1000011001;
    16'b0010000010000001: out_v[111] = 10'b1010101101;
    16'b0010000000000001: out_v[111] = 10'b1001011101;
    16'b0000000010000100: out_v[111] = 10'b1100010101;
    default: out_v[111] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000001000001000: out_v[112] = 10'b1010110001;
    16'b0000100000001000: out_v[112] = 10'b1010100101;
    16'b0000101000000000: out_v[112] = 10'b0111001010;
    16'b0000000000001000: out_v[112] = 10'b1000110111;
    16'b0000001000000000: out_v[112] = 10'b0000001011;
    16'b0000100000000000: out_v[112] = 10'b1100000110;
    16'b0000000000000000: out_v[112] = 10'b0101000111;
    16'b0000101000001000: out_v[112] = 10'b1010111001;
    16'b0000000001001000: out_v[112] = 10'b1000001111;
    16'b0000001001001000: out_v[112] = 10'b0110110001;
    16'b0000000000101000: out_v[112] = 10'b0101110100;
    16'b0000000000100000: out_v[112] = 10'b0000101100;
    16'b0000100000100000: out_v[112] = 10'b0011000110;
    16'b0000001001000000: out_v[112] = 10'b1100100000;
    16'b0000101001001000: out_v[112] = 10'b0101001100;
    16'b0000100001001000: out_v[112] = 10'b0101011100;
    16'b0000100000101000: out_v[112] = 10'b1100011100;
    16'b0000000001000000: out_v[112] = 10'b1111100111;
    16'b0000100001000000: out_v[112] = 10'b1101100111;
    16'b0000101001000000: out_v[112] = 10'b1001110010;
    16'b0000100001100000: out_v[112] = 10'b0011100100;
    16'b0000100001101000: out_v[112] = 10'b0111000000;
    16'b0000000001100000: out_v[112] = 10'b0100100101;
    16'b0000100001101001: out_v[112] = 10'b0000000111;
    16'b0000000001101000: out_v[112] = 10'b0101000110;
    16'b0001100001101000: out_v[112] = 10'b1011011011;
    16'b0000000001101001: out_v[112] = 10'b1101010011;
    16'b0001000001001000: out_v[112] = 10'b1011001010;
    16'b0001100000001000: out_v[112] = 10'b1010100111;
    16'b0000100001100001: out_v[112] = 10'b0111000010;
    16'b0001000000000000: out_v[112] = 10'b1011010010;
    16'b0110000001001000: out_v[112] = 10'b0000001001;
    16'b0001001001000000: out_v[112] = 10'b0100111011;
    16'b0001100001001000: out_v[112] = 10'b1101001001;
    16'b0001000001000000: out_v[112] = 10'b1101100101;
    16'b0001001001001000: out_v[112] = 10'b0011010010;
    16'b0010001001001000: out_v[112] = 10'b0011111110;
    16'b0110001001001000: out_v[112] = 10'b1100110110;
    16'b0001000000001000: out_v[112] = 10'b0000110111;
    16'b0110001000001000: out_v[112] = 10'b0111100000;
    16'b0110000000000000: out_v[112] = 10'b0100100100;
    16'b0110001000000000: out_v[112] = 10'b0011101011;
    16'b0010000001001000: out_v[112] = 10'b1001110001;
    16'b0000001100001000: out_v[112] = 10'b0101110110;
    16'b0110000000001000: out_v[112] = 10'b0110111011;
    16'b0000000101001000: out_v[112] = 10'b1010011000;
    16'b0010000000001000: out_v[112] = 10'b0011110000;
    16'b0000000100001000: out_v[112] = 10'b0110111000;
    16'b0100000001001000: out_v[112] = 10'b1011110001;
    16'b0000001101001000: out_v[112] = 10'b0011011100;
    16'b0010001000001000: out_v[112] = 10'b1101101110;
    16'b0100010001001000: out_v[112] = 10'b1100111011;
    16'b0110000001000000: out_v[112] = 10'b0101101000;
    16'b0100001001001000: out_v[112] = 10'b0101110100;
    16'b0110001001000000: out_v[112] = 10'b1000100111;
    default: out_v[112] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000100100000000: out_v[113] = 10'b0000110011;
    16'b0000100100000010: out_v[113] = 10'b1000101010;
    16'b0000110100001000: out_v[113] = 10'b0101010111;
    16'b0000100101001010: out_v[113] = 10'b1011111010;
    16'b0000100101000000: out_v[113] = 10'b1110010001;
    16'b0000100001000000: out_v[113] = 10'b1001101001;
    16'b0000100000001000: out_v[113] = 10'b1000111011;
    16'b0000000000001000: out_v[113] = 10'b1100100001;
    16'b0000000101001000: out_v[113] = 10'b0100011001;
    16'b0000000100000000: out_v[113] = 10'b0010110010;
    16'b0000100101000010: out_v[113] = 10'b0001011111;
    16'b0010100101000000: out_v[113] = 10'b0110001111;
    16'b0000110100000000: out_v[113] = 10'b1001110000;
    16'b0000100000000000: out_v[113] = 10'b0010000101;
    16'b0000110110001000: out_v[113] = 10'b1111010011;
    16'b0000100110000000: out_v[113] = 10'b1101110001;
    16'b0000100101001000: out_v[113] = 10'b0011110111;
    16'b0000100100001010: out_v[113] = 10'b1011001111;
    16'b0000100001000010: out_v[113] = 10'b0011011110;
    16'b0000110110101000: out_v[113] = 10'b1111000111;
    16'b0000000000000000: out_v[113] = 10'b1000100010;
    16'b0000100000000010: out_v[113] = 10'b1010000111;
    16'b0000100111000000: out_v[113] = 10'b1010100010;
    16'b0000010100101000: out_v[113] = 10'b1010010011;
    16'b0000000100001000: out_v[113] = 10'b0101110111;
    16'b0000100100001000: out_v[113] = 10'b0111101111;
    16'b0000000001001000: out_v[113] = 10'b0001101100;
    16'b0000000100001010: out_v[113] = 10'b1111001111;
    16'b0000100000001010: out_v[113] = 10'b0001110011;
    16'b0000110100101000: out_v[113] = 10'b0000110101;
    16'b0010100100000000: out_v[113] = 10'b1000001100;
    16'b0000010100001000: out_v[113] = 10'b0111011110;
    16'b0000110110000000: out_v[113] = 10'b0111011001;
    16'b0000110100100000: out_v[113] = 10'b0010110110;
    16'b0000100010000000: out_v[113] = 10'b0101001011;
    16'b0010000100000000: out_v[113] = 10'b0101100111;
    16'b0000100001001000: out_v[113] = 10'b1110100111;
    16'b0000000100000010: out_v[113] = 10'b0101000111;
    16'b0000100001001010: out_v[113] = 10'b1110010110;
    16'b0000000101000000: out_v[113] = 10'b0111011100;
    16'b0000110110100000: out_v[113] = 10'b0100001101;
    16'b0000000100101000: out_v[113] = 10'b0011100111;
    16'b0010000000000010: out_v[113] = 10'b1011111011;
    16'b0010000000000000: out_v[113] = 10'b1001101101;
    16'b0010000001000000: out_v[113] = 10'b1101010101;
    16'b0000000010000000: out_v[113] = 10'b0100110110;
    16'b0010000101000000: out_v[113] = 10'b1101000010;
    16'b0010000010000000: out_v[113] = 10'b0011010110;
    16'b0010000110000000: out_v[113] = 10'b1100101110;
    16'b0000000110000000: out_v[113] = 10'b0101001000;
    16'b0010010010000000: out_v[113] = 10'b1001010110;
    16'b0010010010100000: out_v[113] = 10'b0110100001;
    16'b0010010110100000: out_v[113] = 10'b1011100111;
    16'b0010010000000000: out_v[113] = 10'b0011111101;
    16'b0010010011100000: out_v[113] = 10'b1101000011;
    16'b0010000011000000: out_v[113] = 10'b1000111101;
    16'b0010010011000000: out_v[113] = 10'b1000110110;
    16'b0010010110000000: out_v[113] = 10'b0100000101;
    16'b0010100000001000: out_v[113] = 10'b1101001111;
    16'b0000000011000000: out_v[113] = 10'b0100100101;
    16'b0010110011000000: out_v[113] = 10'b1111000011;
    16'b0010100001001000: out_v[113] = 10'b1011001110;
    16'b0010100000000000: out_v[113] = 10'b0101111010;
    16'b0010010111100000: out_v[113] = 10'b1010111001;
    16'b0010000011001000: out_v[113] = 10'b1010011101;
    16'b0010110000000000: out_v[113] = 10'b1001001110;
    16'b0010100001000010: out_v[113] = 10'b0100010001;
    16'b0010010010110000: out_v[113] = 10'b0101111011;
    16'b0010000000001000: out_v[113] = 10'b0100100101;
    16'b0000010010000000: out_v[113] = 10'b0111110100;
    16'b0010000001001000: out_v[113] = 10'b1100101111;
    16'b0010000010100000: out_v[113] = 10'b0111001101;
    16'b0010100001000000: out_v[113] = 10'b0001101001;
    16'b0010100001101000: out_v[113] = 10'b0000100101;
    16'b0000010010100000: out_v[113] = 10'b1011110011;
    16'b0010110010000000: out_v[113] = 10'b0011010011;
    16'b0010100011000000: out_v[113] = 10'b0101010011;
    16'b0010100011001000: out_v[113] = 10'b0110100010;
    16'b0010000011100000: out_v[113] = 10'b1111101100;
    16'b0000000001000000: out_v[113] = 10'b0000110010;
    16'b0010000000100000: out_v[113] = 10'b1000101100;
    16'b0010010000100000: out_v[113] = 10'b0100110111;
    16'b0000010000000000: out_v[113] = 10'b1111001110;
    16'b0010000001100000: out_v[113] = 10'b1001101000;
    16'b0010010100000000: out_v[113] = 10'b1001101010;
    16'b0010110011100000: out_v[113] = 10'b0111001100;
    16'b0010000001000010: out_v[113] = 10'b1110010111;
    16'b0000010100000010: out_v[113] = 10'b0100010111;
    16'b0000010100100000: out_v[113] = 10'b1000001111;
    16'b0000010100000000: out_v[113] = 10'b1010101101;
    16'b0000000000000010: out_v[113] = 10'b0010101111;
    16'b0000010111000010: out_v[113] = 10'b1101010111;
    16'b0000010110000000: out_v[113] = 10'b1001001100;
    16'b0000000111000010: out_v[113] = 10'b1111000101;
    16'b0010010100000010: out_v[113] = 10'b1011001001;
    16'b0010010100100000: out_v[113] = 10'b0010100011;
    16'b0010000100000010: out_v[113] = 10'b0001001010;
    16'b0010110100000000: out_v[113] = 10'b1010100111;
    16'b0000000001000010: out_v[113] = 10'b1011000100;
    16'b0000010111000000: out_v[113] = 10'b0001111011;
    16'b0000000101000010: out_v[113] = 10'b1011011101;
    16'b0000000111000000: out_v[113] = 10'b0010111001;
    16'b0000110100000010: out_v[113] = 10'b1100011110;
    16'b0000010110100000: out_v[113] = 10'b0101110000;
    16'b0010110100000010: out_v[113] = 10'b0111100011;
    16'b0000110111000000: out_v[113] = 10'b0111110010;
    16'b0010000100001000: out_v[113] = 10'b1110110001;
    16'b0010110000001000: out_v[113] = 10'b0110111011;
    16'b0010100100001000: out_v[113] = 10'b1001010100;
    16'b0010100000101000: out_v[113] = 10'b1000110100;
    16'b0000110000000000: out_v[113] = 10'b0000111100;
    16'b0010110000101000: out_v[113] = 10'b1010011110;
    16'b0010110100001000: out_v[113] = 10'b1110011011;
    16'b0010100010000000: out_v[113] = 10'b0111111010;
    16'b0000110010000000: out_v[113] = 10'b1100011101;
    16'b0000001000000000: out_v[113] = 10'b0011010011;
    16'b0000001100000000: out_v[113] = 10'b1010100011;
    16'b0000101100000000: out_v[113] = 10'b0011010001;
    16'b1000101000000000: out_v[113] = 10'b1100111001;
    16'b0000101000000000: out_v[113] = 10'b0010011111;
    16'b1000000000000000: out_v[113] = 10'b1010100111;
    16'b1000001000000000: out_v[113] = 10'b1101011110;
    16'b0010100000000010: out_v[113] = 10'b1000010111;
    16'b0010010111000000: out_v[113] = 10'b1000111011;
    16'b0010100100000010: out_v[113] = 10'b0101100000;
    16'b0010110100100000: out_v[113] = 10'b0110100010;
    16'b0010000111000000: out_v[113] = 10'b1011000011;
    default: out_v[113] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100000000000001: out_v[114] = 10'b0011101011;
    16'b0100000000000101: out_v[114] = 10'b1000110100;
    16'b1000000000000101: out_v[114] = 10'b0101001011;
    16'b0000000000000101: out_v[114] = 10'b0101011001;
    16'b1100000000000100: out_v[114] = 10'b1101011000;
    16'b0000001000000100: out_v[114] = 10'b0011100011;
    16'b0100000000000100: out_v[114] = 10'b0000101010;
    16'b0100001000000100: out_v[114] = 10'b1011101001;
    16'b0000001000000101: out_v[114] = 10'b1000001001;
    16'b0100000000010101: out_v[114] = 10'b0110101100;
    16'b1100000000000101: out_v[114] = 10'b0011111010;
    16'b0000000000000001: out_v[114] = 10'b0010100110;
    16'b0100000000000000: out_v[114] = 10'b0000101111;
    16'b1100000000000001: out_v[114] = 10'b0111000000;
    16'b0100001000000101: out_v[114] = 10'b0001111111;
    16'b1100001000000101: out_v[114] = 10'b1010110111;
    16'b0000001000000001: out_v[114] = 10'b1001000111;
    16'b0000000000000100: out_v[114] = 10'b0010011010;
    16'b1100000000000000: out_v[114] = 10'b1001011000;
    16'b0000000000000000: out_v[114] = 10'b0111010100;
    16'b1000000000000100: out_v[114] = 10'b0011000011;
    16'b1000001000000101: out_v[114] = 10'b0000001011;
    16'b1100000000010001: out_v[114] = 10'b1100010010;
    16'b0000000000010001: out_v[114] = 10'b0011001110;
    16'b0000000000010000: out_v[114] = 10'b1001001100;
    16'b0100000000010001: out_v[114] = 10'b1100000000;
    16'b0100000000010000: out_v[114] = 10'b0001110011;
    16'b1000000000010001: out_v[114] = 10'b1001111110;
    16'b1000000000010000: out_v[114] = 10'b1010100110;
    16'b1100000000010000: out_v[114] = 10'b0101001101;
    16'b0000001000010000: out_v[114] = 10'b0001101111;
    16'b1000001000010000: out_v[114] = 10'b1100101110;
    16'b0000000000011000: out_v[114] = 10'b0011001100;
    16'b0000000000001000: out_v[114] = 10'b1110101110;
    16'b0000001000000000: out_v[114] = 10'b1100010110;
    16'b1000000000000000: out_v[114] = 10'b1100100100;
    16'b0000001000010001: out_v[114] = 10'b0011001110;
    16'b0000001000010100: out_v[114] = 10'b0101110000;
    16'b0000000000010100: out_v[114] = 10'b1101010010;
    16'b1000000000010100: out_v[114] = 10'b1111110101;
    16'b0100001000011000: out_v[114] = 10'b0010100101;
    16'b0100001000010000: out_v[114] = 10'b1000000111;
    16'b0100001000000000: out_v[114] = 10'b0101110010;
    16'b0000000000010101: out_v[114] = 10'b1100010000;
    16'b1000000000000001: out_v[114] = 10'b1011010111;
    16'b0000001000011000: out_v[114] = 10'b1111110111;
    16'b0000000010010001: out_v[114] = 10'b0010101001;
    16'b0100001000010101: out_v[114] = 10'b0110010011;
    16'b0100001000010001: out_v[114] = 10'b1010011001;
    16'b0100000000010100: out_v[114] = 10'b1000010110;
    16'b1100000000010101: out_v[114] = 10'b1000001111;
    16'b0100000010010001: out_v[114] = 10'b0001111000;
    16'b1000000000010101: out_v[114] = 10'b0110110110;
    16'b0100000010010101: out_v[114] = 10'b0101101001;
    16'b0000000010010101: out_v[114] = 10'b1100100101;
    16'b0000000001010100: out_v[114] = 10'b0010010111;
    16'b0100000010000101: out_v[114] = 10'b0101110010;
    16'b0100000010000001: out_v[114] = 10'b0101111110;
    16'b0000001000010101: out_v[114] = 10'b1100010010;
    16'b1100000000010100: out_v[114] = 10'b0111011100;
    16'b0000001000011100: out_v[114] = 10'b1111000110;
    16'b0000000000011100: out_v[114] = 10'b1001001010;
    16'b1101000000000000: out_v[114] = 10'b1001011010;
    16'b1000001000010100: out_v[114] = 10'b1001010010;
    16'b1101000000010100: out_v[114] = 10'b1100010101;
    16'b1101000000010000: out_v[114] = 10'b1110111101;
    16'b0100001000010100: out_v[114] = 10'b0110110010;
    16'b0000000010000101: out_v[114] = 10'b0011010111;
    16'b0000000010000001: out_v[114] = 10'b0010110000;
    16'b0000000010010000: out_v[114] = 10'b0110011001;
    16'b0100000001000100: out_v[114] = 10'b1110001110;
    16'b0000000010010100: out_v[114] = 10'b1101010011;
    16'b0000000010000000: out_v[114] = 10'b1100001011;
    16'b0100000010010100: out_v[114] = 10'b0101011011;
    16'b0100000010010000: out_v[114] = 10'b1100001110;
    16'b0000000001000000: out_v[114] = 10'b1001010011;
    default: out_v[114] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010100001100000: out_v[115] = 10'b1001010101;
    16'b0011100001100000: out_v[115] = 10'b1101001110;
    16'b0011100001000000: out_v[115] = 10'b0111100001;
    16'b0011100001101000: out_v[115] = 10'b1100100101;
    16'b0000000001100000: out_v[115] = 10'b1000001111;
    16'b0010100000000000: out_v[115] = 10'b0000100001;
    16'b0001100000001000: out_v[115] = 10'b1011010111;
    16'b0001000000101000: out_v[115] = 10'b1010010111;
    16'b0000100001000000: out_v[115] = 10'b1100100101;
    16'b0001000000000000: out_v[115] = 10'b0100011001;
    16'b0001100000101000: out_v[115] = 10'b1000111101;
    16'b0001100001001000: out_v[115] = 10'b1001011111;
    16'b0001100000100000: out_v[115] = 10'b0110011111;
    16'b0001100001100000: out_v[115] = 10'b1001010011;
    16'b0010100001000000: out_v[115] = 10'b0111011001;
    16'b0001000000100000: out_v[115] = 10'b1100001111;
    16'b0011100001001000: out_v[115] = 10'b1001010111;
    16'b0000000001000000: out_v[115] = 10'b0100001101;
    16'b0010100001101000: out_v[115] = 10'b0111001111;
    16'b0000100001100000: out_v[115] = 10'b0100010111;
    16'b0001100001000000: out_v[115] = 10'b0110100110;
    16'b0001000001100000: out_v[115] = 10'b1110111011;
    16'b0001100001101000: out_v[115] = 10'b0010111110;
    16'b0010000001000000: out_v[115] = 10'b0100001110;
    16'b0010100000100000: out_v[115] = 10'b1000110101;
    16'b0010000001100000: out_v[115] = 10'b1000011111;
    16'b0001100000000000: out_v[115] = 10'b1100011111;
    16'b0010000000000000: out_v[115] = 10'b1010100010;
    16'b0000100001101000: out_v[115] = 10'b0111011011;
    16'b0001000001000000: out_v[115] = 10'b1010111010;
    16'b0010100001001000: out_v[115] = 10'b1111010001;
    16'b0000100000100000: out_v[115] = 10'b0111001000;
    16'b0010001001100000: out_v[115] = 10'b0100011000;
    16'b0010101001100000: out_v[115] = 10'b1100001110;
    16'b0000101000000000: out_v[115] = 10'b0111011110;
    16'b0000101000100000: out_v[115] = 10'b0010100000;
    16'b0010101000100000: out_v[115] = 10'b1000100010;
    16'b0010001001000000: out_v[115] = 10'b0000011010;
    16'b0000001000000000: out_v[115] = 10'b0011100100;
    16'b0010001000100000: out_v[115] = 10'b0101111101;
    16'b0000100000000000: out_v[115] = 10'b0101011110;
    16'b0000001000100000: out_v[115] = 10'b0011110001;
    16'b0010101001000000: out_v[115] = 10'b1110001000;
    16'b0010101000000000: out_v[115] = 10'b1101100000;
    16'b0010001000000000: out_v[115] = 10'b0111000000;
    16'b0011001001000000: out_v[115] = 10'b1001010110;
    16'b0000000000000000: out_v[115] = 10'b0001101010;
    16'b0000111010000000: out_v[115] = 10'b1010000111;
    16'b0010111000000000: out_v[115] = 10'b1111100100;
    16'b0010001001101000: out_v[115] = 10'b0000011111;
    16'b0010011001100000: out_v[115] = 10'b1110010101;
    16'b0010101001101000: out_v[115] = 10'b1011011101;
    16'b0010000001101000: out_v[115] = 10'b1000001010;
    16'b0010010011100000: out_v[115] = 10'b0101001101;
    16'b0010011011100000: out_v[115] = 10'b0100011000;
    16'b0010101001001000: out_v[115] = 10'b0011011011;
    16'b0010110010000000: out_v[115] = 10'b1100010111;
    16'b0010111010000000: out_v[115] = 10'b1010001000;
    16'b0000111000000000: out_v[115] = 10'b1111001010;
    16'b0010000001001000: out_v[115] = 10'b0110010001;
    16'b0010101000001000: out_v[115] = 10'b0011001001;
    16'b0010001001001000: out_v[115] = 10'b1110000111;
    16'b0000111010010000: out_v[115] = 10'b0101011000;
    16'b0011101000101000: out_v[115] = 10'b1111011010;
    16'b0011101001101000: out_v[115] = 10'b1110101011;
    16'b0011101001000000: out_v[115] = 10'b1010101100;
    16'b0011001000101000: out_v[115] = 10'b0010011000;
    16'b0011101001001000: out_v[115] = 10'b0001110100;
    16'b0011001001101000: out_v[115] = 10'b1001010100;
    16'b0000101000010000: out_v[115] = 10'b0010110101;
    16'b0011001000000000: out_v[115] = 10'b0011110010;
    16'b0001001000000000: out_v[115] = 10'b0100011011;
    16'b0010001001010000: out_v[115] = 10'b0000011111;
    16'b0011000000000000: out_v[115] = 10'b0001110000;
    16'b0010000000010000: out_v[115] = 10'b0111010110;
    16'b0011101000000000: out_v[115] = 10'b0100010011;
    16'b0010101000010000: out_v[115] = 10'b1101100010;
    16'b0010000000100000: out_v[115] = 10'b0000110111;
    16'b0010001000010000: out_v[115] = 10'b0011001110;
    16'b0010000001010000: out_v[115] = 10'b1001011010;
    16'b0011100000000000: out_v[115] = 10'b0011111100;
    16'b0011000001000000: out_v[115] = 10'b1001100000;
    16'b0001101001000000: out_v[115] = 10'b1000100110;
    16'b0000101001000000: out_v[115] = 10'b1100100011;
    16'b0001101001100000: out_v[115] = 10'b1001101110;
    16'b0000101000101000: out_v[115] = 10'b1101111001;
    16'b0001101001001000: out_v[115] = 10'b0110001010;
    16'b0001101000000000: out_v[115] = 10'b0100011111;
    16'b0000000000100000: out_v[115] = 10'b1010100000;
    16'b0000101000001000: out_v[115] = 10'b1111110010;
    16'b0000001000101000: out_v[115] = 10'b0001110111;
    16'b0011100101000000: out_v[115] = 10'b0110011100;
    16'b0010100101000000: out_v[115] = 10'b0111111001;
    16'b0010101101000000: out_v[115] = 10'b1000101101;
    16'b0010100000010000: out_v[115] = 10'b1101100011;
    16'b0011100100000000: out_v[115] = 10'b1111111100;
    16'b0010100100000000: out_v[115] = 10'b1011100010;
    16'b0001100101000000: out_v[115] = 10'b0011010111;
    16'b0010101100000000: out_v[115] = 10'b1001100101;
    16'b0011101101000000: out_v[115] = 10'b1101000100;
    16'b0011101001100000: out_v[115] = 10'b0111100110;
    16'b0001101000100000: out_v[115] = 10'b0001011011;
    16'b0011101000100000: out_v[115] = 10'b0110011100;
    16'b0001001000100000: out_v[115] = 10'b1110001010;
    16'b0011001000100000: out_v[115] = 10'b0001001010;
    16'b0011001001100000: out_v[115] = 10'b1110000001;
    16'b0010101001010000: out_v[115] = 10'b1001100101;
    16'b0010100001010000: out_v[115] = 10'b1000101110;
    16'b0010111010010000: out_v[115] = 10'b0110000101;
    default: out_v[115] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000001000010001: out_v[116] = 10'b0010101111;
    16'b0000011010001011: out_v[116] = 10'b1010100011;
    16'b1010000000001111: out_v[116] = 10'b0111111111;
    16'b0010000000011001: out_v[116] = 10'b0011001011;
    16'b0000000000001001: out_v[116] = 10'b1101110111;
    16'b1000001000000101: out_v[116] = 10'b0010100111;
    16'b1010010010001111: out_v[116] = 10'b1111110011;
    16'b1000000000001001: out_v[116] = 10'b0100110011;
    16'b0000000000010001: out_v[116] = 10'b1101010001;
    16'b0010001000011001: out_v[116] = 10'b1110110111;
    16'b1000011010001111: out_v[116] = 10'b1010101101;
    16'b1000000000011001: out_v[116] = 10'b0001011110;
    16'b1000000000000101: out_v[116] = 10'b0011001000;
    16'b1000001000001101: out_v[116] = 10'b1111001111;
    16'b0000000000000001: out_v[116] = 10'b1101100001;
    16'b1000000000001100: out_v[116] = 10'b1101011001;
    16'b0000000000011001: out_v[116] = 10'b1000111000;
    16'b1000000000001111: out_v[116] = 10'b1110111010;
    16'b1000010010001101: out_v[116] = 10'b0111011011;
    16'b1010000000001101: out_v[116] = 10'b1110011010;
    16'b1010000000010001: out_v[116] = 10'b0010110010;
    16'b1000000000001101: out_v[116] = 10'b1001111110;
    16'b1000000000000100: out_v[116] = 10'b1110011011;
    16'b0000011010011011: out_v[116] = 10'b1010111111;
    16'b1010000000001001: out_v[116] = 10'b0000111111;
    16'b1000000000010001: out_v[116] = 10'b0100101110;
    16'b0000011010001111: out_v[116] = 10'b0111011011;
    16'b1000010010001111: out_v[116] = 10'b1101010011;
    16'b1000001000001111: out_v[116] = 10'b0111011111;
    16'b0000001000011001: out_v[116] = 10'b1110100100;
    16'b1000001000011101: out_v[116] = 10'b1101001000;
    16'b0010001000010001: out_v[116] = 10'b0011011000;
    16'b0000001000011011: out_v[116] = 10'b0010001101;
    16'b1000000000000001: out_v[116] = 10'b0010110101;
    16'b1000000000000000: out_v[116] = 10'b1000101001;
    16'b0010000000001001: out_v[116] = 10'b0111000110;
    16'b1000000000011101: out_v[116] = 10'b1100011110;
    16'b1000001000010001: out_v[116] = 10'b1101100110;
    16'b1010000000011001: out_v[116] = 10'b1011000110;
    16'b0010000000010001: out_v[116] = 10'b1011011010;
    16'b1000000100001100: out_v[116] = 10'b0111100110;
    16'b0010000000000001: out_v[116] = 10'b1101110001;
    16'b1010000000001100: out_v[116] = 10'b1110111011;
    16'b1010000000000001: out_v[116] = 10'b1010110100;
    16'b0000011010011001: out_v[116] = 10'b1010110101;
    16'b0000001000001111: out_v[116] = 10'b1001100011;
    16'b1000001000011001: out_v[116] = 10'b0101110111;
    16'b0000010010011000: out_v[116] = 10'b1010100101;
    16'b0000000000001000: out_v[116] = 10'b0011111010;
    16'b0000001000000000: out_v[116] = 10'b0011001010;
    16'b0000000000000000: out_v[116] = 10'b0111101001;
    16'b0000001000010000: out_v[116] = 10'b0101110011;
    16'b0000000000011000: out_v[116] = 10'b0011111101;
    16'b0000001000000001: out_v[116] = 10'b1111001011;
    16'b0000000000010000: out_v[116] = 10'b0010101100;
    16'b0010001000000000: out_v[116] = 10'b1101100010;
    16'b0000001000011000: out_v[116] = 10'b1111110001;
    16'b0000010000011010: out_v[116] = 10'b1111110011;
    16'b0000010010011010: out_v[116] = 10'b1010110111;
    16'b0010001000010000: out_v[116] = 10'b1111110010;
    16'b0000010000011000: out_v[116] = 10'b1011111011;
    16'b0001010010011010: out_v[116] = 10'b0001011111;
    16'b0000001000001000: out_v[116] = 10'b0101110001;
    16'b0010000000000000: out_v[116] = 10'b1101101010;
    16'b0000011010011000: out_v[116] = 10'b1111000001;
    16'b0000011000011000: out_v[116] = 10'b0011101010;
    16'b0000010000001000: out_v[116] = 10'b1111101101;
    16'b0010000000010000: out_v[116] = 10'b1100100100;
    16'b0010000000010010: out_v[116] = 10'b1000100100;
    16'b0010000000011000: out_v[116] = 10'b1000100110;
    16'b0000000000000100: out_v[116] = 10'b1010100111;
    16'b0010000000000010: out_v[116] = 10'b1100100110;
    16'b0010000000001010: out_v[116] = 10'b1011011000;
    16'b0010000000011010: out_v[116] = 10'b1000110100;
    16'b0010000000011100: out_v[116] = 10'b1111101010;
    16'b0010000000011110: out_v[116] = 10'b1011011011;
    16'b0000000000011010: out_v[116] = 10'b1011011110;
    16'b0010000000010100: out_v[116] = 10'b1110100101;
    16'b0000000000010100: out_v[116] = 10'b0011100110;
    16'b0000000100000000: out_v[116] = 10'b1101100100;
    16'b0000000100010000: out_v[116] = 10'b1011111010;
    16'b0010010010011010: out_v[116] = 10'b1010110100;
    16'b0010000000001100: out_v[116] = 10'b1010011011;
    16'b0000000000010010: out_v[116] = 10'b1001101110;
    16'b0000001000110000: out_v[116] = 10'b0010000101;
    16'b0000010010011100: out_v[116] = 10'b1010101110;
    16'b0010010010011110: out_v[116] = 10'b0111111001;
    16'b0000001000010100: out_v[116] = 10'b1000100110;
    16'b0010010000011010: out_v[116] = 10'b1111010101;
    16'b0000000000110000: out_v[116] = 10'b1101000110;
    16'b0000000000011100: out_v[116] = 10'b0110100111;
    16'b0000001000000010: out_v[116] = 10'b1101111000;
    16'b0000000000000010: out_v[116] = 10'b0000111111;
    16'b0000000000001010: out_v[116] = 10'b1000011010;
    16'b0000001100000000: out_v[116] = 10'b1000001110;
    16'b0010010010001010: out_v[116] = 10'b1010100100;
    16'b0010001000000011: out_v[116] = 10'b1111010100;
    16'b0000010010001010: out_v[116] = 10'b1001011011;
    16'b0000001000001010: out_v[116] = 10'b0010010100;
    16'b1000001000000001: out_v[116] = 10'b1010001000;
    16'b0001000000001010: out_v[116] = 10'b0010110011;
    16'b0010001000000010: out_v[116] = 10'b0111010001;
    16'b0010001000000001: out_v[116] = 10'b0100011111;
    16'b0010000000001000: out_v[116] = 10'b1001111100;
    16'b0000001000001011: out_v[116] = 10'b0011101111;
    16'b0000001000000011: out_v[116] = 10'b0000011110;
    16'b0001000000000010: out_v[116] = 10'b0010100000;
    16'b0001010010001010: out_v[116] = 10'b0001011110;
    16'b0010001000001010: out_v[116] = 10'b1011011011;
    16'b0010001000001011: out_v[116] = 10'b0010011110;
    16'b0001001000001010: out_v[116] = 10'b1001010100;
    16'b1000000000011000: out_v[116] = 10'b0111010011;
    16'b1000010010001001: out_v[116] = 10'b1001011000;
    16'b1000000000011100: out_v[116] = 10'b1101111011;
    16'b0000010010001001: out_v[116] = 10'b1110101001;
    16'b0000010010011001: out_v[116] = 10'b1010110110;
    16'b0000010000011001: out_v[116] = 10'b1111011000;
    16'b1000010010011101: out_v[116] = 10'b0111110000;
    16'b0000000000011101: out_v[116] = 10'b0111110110;
    16'b1000000000001000: out_v[116] = 10'b1101100100;
    16'b1000010010011001: out_v[116] = 10'b0110101111;
    16'b1000000000010000: out_v[116] = 10'b1101010010;
    16'b0000010010011101: out_v[116] = 10'b1110110010;
    16'b0000000000010101: out_v[116] = 10'b1101011000;
    16'b1000000000010101: out_v[116] = 10'b0000110010;
    16'b1000000000010100: out_v[116] = 10'b1101011000;
    16'b1000010010011100: out_v[116] = 10'b0110100011;
    16'b0000010000001001: out_v[116] = 10'b1110010111;
    16'b1000000010001001: out_v[116] = 10'b0110111110;
    16'b0000001000010101: out_v[116] = 10'b0000011011;
    16'b1000000010011001: out_v[116] = 10'b1001100011;
    16'b0000000000000101: out_v[116] = 10'b0100110010;
    16'b0000010010001101: out_v[116] = 10'b1110101010;
    16'b0000001000001001: out_v[116] = 10'b0111110110;
    16'b0000011010001001: out_v[116] = 10'b0010110110;
    16'b0000000010001001: out_v[116] = 10'b0010111101;
    16'b1000010010001011: out_v[116] = 10'b1001111010;
    16'b0000011010001000: out_v[116] = 10'b1000110111;
    16'b0000011010001010: out_v[116] = 10'b1010111111;
    16'b0000010000000001: out_v[116] = 10'b0010111010;
    16'b0000010010001011: out_v[116] = 10'b1010101011;
    16'b0000001010001001: out_v[116] = 10'b0011111101;
    16'b1000011010001001: out_v[116] = 10'b1010101100;
    16'b1000001000001001: out_v[116] = 10'b1111100001;
    16'b1000011010001011: out_v[116] = 10'b1000100110;
    16'b0000000000001011: out_v[116] = 10'b1001110011;
    16'b1000001000001011: out_v[116] = 10'b1111111010;
    16'b0000011000010000: out_v[116] = 10'b1011011010;
    16'b1010000000000101: out_v[116] = 10'b1101011111;
    16'b1000000000110001: out_v[116] = 10'b0111011100;
    16'b1000000000110000: out_v[116] = 10'b0011111011;
    16'b1010000000010101: out_v[116] = 10'b0111110010;
    16'b0000011000010001: out_v[116] = 10'b1001011110;
    16'b1000001100000001: out_v[116] = 10'b0010110001;
    16'b0000001100000001: out_v[116] = 10'b1010011000;
    16'b0000000100001000: out_v[116] = 10'b1001110011;
    16'b1000000100000001: out_v[116] = 10'b0111100010;
    16'b1000001100000000: out_v[116] = 10'b1011001001;
    16'b0000001001001001: out_v[116] = 10'b1101101001;
    16'b1000001000000000: out_v[116] = 10'b1001000111;
    16'b1000001001001001: out_v[116] = 10'b0011111000;
    16'b1000000001001001: out_v[116] = 10'b1110111011;
    16'b1000000100000000: out_v[116] = 10'b1001011111;
    16'b1000001100001001: out_v[116] = 10'b0111100000;
    16'b0000000001001000: out_v[116] = 10'b0111011010;
    16'b1000001001000001: out_v[116] = 10'b0111010110;
    16'b0000000000011011: out_v[116] = 10'b0111110110;
    16'b0000011010011010: out_v[116] = 10'b1000100101;
    16'b0001010010011011: out_v[116] = 10'b0101010000;
    16'b0000001000011010: out_v[116] = 10'b1101110001;
    16'b0001011010011010: out_v[116] = 10'b0100100010;
    16'b0000010010011011: out_v[116] = 10'b1111010011;
    16'b1000000100010001: out_v[116] = 10'b1111000010;
    16'b0000000010011001: out_v[116] = 10'b0100111010;
    16'b0010001000011000: out_v[116] = 10'b1100000011;
    16'b1000010010011011: out_v[116] = 10'b1100000100;
    16'b1000000100010100: out_v[116] = 10'b1101111110;
    16'b1000000100010000: out_v[116] = 10'b0001010001;
    default: out_v[116] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0101100010010000: out_v[117] = 10'b0111001011;
    16'b0101100010011000: out_v[117] = 10'b1000100011;
    16'b0001101010011000: out_v[117] = 10'b0001100101;
    16'b0101100000001000: out_v[117] = 10'b0100010111;
    16'b0101100010000000: out_v[117] = 10'b1000101001;
    16'b0001100000011000: out_v[117] = 10'b0001001001;
    16'b0001001010001000: out_v[117] = 10'b1001010010;
    16'b0100100000011000: out_v[117] = 10'b0000000100;
    16'b0101001010001000: out_v[117] = 10'b1001001111;
    16'b0001000010001000: out_v[117] = 10'b1001101010;
    16'b0001100010010000: out_v[117] = 10'b1001001010;
    16'b0101101010011000: out_v[117] = 10'b1101010011;
    16'b0101100000011000: out_v[117] = 10'b0101001011;
    16'b0101100010001000: out_v[117] = 10'b0011101001;
    16'b0001101000011000: out_v[117] = 10'b1010001111;
    16'b0001100010011000: out_v[117] = 10'b1001101100;
    16'b0000101010011000: out_v[117] = 10'b0011100011;
    16'b0101101010101000: out_v[117] = 10'b1101100111;
    16'b0101101010111000: out_v[117] = 10'b0000010011;
    16'b0001100010000000: out_v[117] = 10'b0101001001;
    16'b0101101010001000: out_v[117] = 10'b1001101000;
    16'b0000100010011000: out_v[117] = 10'b0011101010;
    16'b0100100010000000: out_v[117] = 10'b0010011010;
    16'b0101100000010000: out_v[117] = 10'b1001110010;
    16'b0100100010011000: out_v[117] = 10'b1001000100;
    16'b0001100010001000: out_v[117] = 10'b1011110000;
    16'b0100000010001000: out_v[117] = 10'b1110001001;
    16'b0101000010001000: out_v[117] = 10'b0110111110;
    16'b0101101000011000: out_v[117] = 10'b1110111011;
    16'b0101100000000000: out_v[117] = 10'b0011001010;
    16'b0100100010010000: out_v[117] = 10'b0001011111;
    16'b0100000010010000: out_v[117] = 10'b0110111011;
    16'b0000100010010000: out_v[117] = 10'b1010011000;
    16'b0000100000000000: out_v[117] = 10'b1011110010;
    16'b0000000000000000: out_v[117] = 10'b1101011111;
    16'b0000000010000000: out_v[117] = 10'b1010111001;
    16'b0000000010010000: out_v[117] = 10'b0011000010;
    16'b0100000010000000: out_v[117] = 10'b0000111111;
    16'b0001000000000000: out_v[117] = 10'b1001101011;
    16'b0000100010000000: out_v[117] = 10'b0110101001;
    16'b0100000010011000: out_v[117] = 10'b0111101011;
    16'b0100000000001000: out_v[117] = 10'b1010101010;
    16'b0000100000010000: out_v[117] = 10'b0110110000;
    16'b0001100000000000: out_v[117] = 10'b1101100110;
    16'b0101000010110000: out_v[117] = 10'b1111110111;
    16'b0101000010010000: out_v[117] = 10'b0101000101;
    16'b0100100000010000: out_v[117] = 10'b1101100001;
    16'b0101100010100000: out_v[117] = 10'b1001110111;
    16'b0101000000010000: out_v[117] = 10'b0001101101;
    16'b0100000010100000: out_v[117] = 10'b0000101111;
    16'b0101000000011000: out_v[117] = 10'b1111010011;
    16'b0101000000001000: out_v[117] = 10'b0001010101;
    16'b0101000010000000: out_v[117] = 10'b1010100110;
    16'b0100000000010000: out_v[117] = 10'b1101000100;
    16'b0101100010110000: out_v[117] = 10'b1010010110;
    16'b0101000000000000: out_v[117] = 10'b1010000011;
    16'b0001000010010000: out_v[117] = 10'b1101011111;
    16'b0001000010000000: out_v[117] = 10'b0001110111;
    16'b0101000000100000: out_v[117] = 10'b0001100010;
    16'b0101000010100000: out_v[117] = 10'b0010011100;
    16'b0001000000001000: out_v[117] = 10'b0100111110;
    16'b0100000000100000: out_v[117] = 10'b1001101111;
    16'b0001000000011000: out_v[117] = 10'b1111001100;
    16'b0100000000000000: out_v[117] = 10'b0000101100;
    16'b0001100000010000: out_v[117] = 10'b0010100010;
    16'b0000000000001000: out_v[117] = 10'b0001111100;
    16'b0101000010011000: out_v[117] = 10'b1100010111;
    16'b0100000000011000: out_v[117] = 10'b0110000001;
    16'b0001100000001000: out_v[117] = 10'b1011111100;
    16'b0000100000011000: out_v[117] = 10'b0000011011;
    16'b0000100000001000: out_v[117] = 10'b0100010111;
    16'b0000101000001000: out_v[117] = 10'b0101011111;
    16'b0100100000001000: out_v[117] = 10'b0101011000;
    16'b0001101000001000: out_v[117] = 10'b0000010110;
    16'b0000000000011000: out_v[117] = 10'b0010011110;
    16'b0100100000000000: out_v[117] = 10'b1111000000;
    16'b0000000000010000: out_v[117] = 10'b1001011001;
    16'b0001001000001000: out_v[117] = 10'b0001110110;
    16'b0001001010000000: out_v[117] = 10'b0101010000;
    16'b0000101010000000: out_v[117] = 10'b0111110101;
    16'b0101001000001000: out_v[117] = 10'b0101001011;
    16'b0001001000000000: out_v[117] = 10'b0011000010;
    16'b0000100010001000: out_v[117] = 10'b1110101011;
    16'b0000000010001000: out_v[117] = 10'b1100101001;
    16'b0000000010011000: out_v[117] = 10'b1111001011;
    16'b0101001000000000: out_v[117] = 10'b1011110010;
    16'b0001101010001000: out_v[117] = 10'b1111000110;
    16'b0001000010001100: out_v[117] = 10'b1110100110;
    16'b0001000000000100: out_v[117] = 10'b1101000111;
    16'b0001000010000100: out_v[117] = 10'b0110000111;
    16'b0000100010000100: out_v[117] = 10'b1101101111;
    16'b0000000010000100: out_v[117] = 10'b1001100100;
    16'b0001100010000100: out_v[117] = 10'b0111110111;
    16'b0000100010001100: out_v[117] = 10'b1011011010;
    16'b0001100010001100: out_v[117] = 10'b0000111110;
    16'b0000000000000100: out_v[117] = 10'b1111101001;
    16'b1000100010000000: out_v[117] = 10'b1000101001;
    16'b0000101010001000: out_v[117] = 10'b1001101011;
    16'b0100100010001000: out_v[117] = 10'b0110010100;
    16'b0101001010000000: out_v[117] = 10'b1000011111;
    16'b0001000010000001: out_v[117] = 10'b1110000101;
    16'b0001000011000000: out_v[117] = 10'b1101101111;
    default: out_v[117] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100010000010010: out_v[118] = 10'b1000011011;
    16'b0100011000000010: out_v[118] = 10'b0010101111;
    16'b0000001100000001: out_v[118] = 10'b0001001111;
    16'b0100001100000000: out_v[118] = 10'b0010010001;
    16'b0000001110000000: out_v[118] = 10'b0010001111;
    16'b0000011000000000: out_v[118] = 10'b1001001011;
    16'b0100001100000001: out_v[118] = 10'b1000101001;
    16'b0000010000010010: out_v[118] = 10'b1011010001;
    16'b0000001100000000: out_v[118] = 10'b0111011101;
    16'b0100011000000000: out_v[118] = 10'b1001110010;
    16'b0100011000000011: out_v[118] = 10'b1110001011;
    16'b0100011100000010: out_v[118] = 10'b0100110001;
    16'b0000011000000010: out_v[118] = 10'b0001011110;
    16'b0000011100000010: out_v[118] = 10'b0011000011;
    16'b0000011100000000: out_v[118] = 10'b1101010110;
    16'b0100011100010000: out_v[118] = 10'b1111100000;
    16'b0100011000010000: out_v[118] = 10'b1111100001;
    16'b0100011000010010: out_v[118] = 10'b1001001000;
    16'b0000011000010010: out_v[118] = 10'b0111101001;
    16'b0000011000000011: out_v[118] = 10'b1111011011;
    16'b0100010000010000: out_v[118] = 10'b1010101111;
    16'b0100010000000010: out_v[118] = 10'b0101010000;
    16'b0100011100010010: out_v[118] = 10'b1001100011;
    16'b0100011100000000: out_v[118] = 10'b1101111100;
    16'b0100001000000000: out_v[118] = 10'b1000011101;
    16'b0100011000000001: out_v[118] = 10'b1110111011;
    16'b0000010000000010: out_v[118] = 10'b1101111001;
    16'b0100011100000011: out_v[118] = 10'b1100001101;
    16'b0000011100000001: out_v[118] = 10'b1111001111;
    16'b0000000110000000: out_v[118] = 10'b0000011101;
    16'b0000001000000000: out_v[118] = 10'b1001000111;
    16'b0000011100010010: out_v[118] = 10'b0100110011;
    16'b0100001100010000: out_v[118] = 10'b0011010001;
    16'b0100010000000000: out_v[118] = 10'b0110100100;
    16'b0100011100000001: out_v[118] = 10'b1011110110;
    16'b0000000100000000: out_v[118] = 10'b0011000101;
    16'b0100001110000000: out_v[118] = 10'b1111010011;
    16'b0100000000000000: out_v[118] = 10'b1100100101;
    16'b0000000000000000: out_v[118] = 10'b1000011011;
    16'b0000010000000000: out_v[118] = 10'b0111001011;
    16'b0100000000000010: out_v[118] = 10'b0001000110;
    16'b0000000000000010: out_v[118] = 10'b0110001011;
    16'b0000000000001000: out_v[118] = 10'b0001010110;
    16'b0000000000010000: out_v[118] = 10'b1100000100;
    16'b0100000000010010: out_v[118] = 10'b1000101110;
    16'b0100000000010000: out_v[118] = 10'b1100001110;
    16'b0000000010000010: out_v[118] = 10'b0110100110;
    16'b0000000000011010: out_v[118] = 10'b0101010111;
    16'b0100001000010000: out_v[118] = 10'b0101110010;
    16'b0100001000010010: out_v[118] = 10'b1000101110;
    16'b0000000000001010: out_v[118] = 10'b1011010111;
    16'b0000001000000010: out_v[118] = 10'b1111000101;
    16'b0100000000011000: out_v[118] = 10'b1110011111;
    16'b0000011010000010: out_v[118] = 10'b0100000111;
    16'b0000001000010010: out_v[118] = 10'b0110000010;
    16'b0000001000010000: out_v[118] = 10'b1111101010;
    16'b0000000000010010: out_v[118] = 10'b1011001111;
    16'b0000001010000000: out_v[118] = 10'b1101001000;
    16'b0000001010010010: out_v[118] = 10'b0001101111;
    16'b0100000000001010: out_v[118] = 10'b0111110011;
    16'b0000000000011000: out_v[118] = 10'b1001100101;
    16'b0100000000011010: out_v[118] = 10'b1011110110;
    16'b0000011010010010: out_v[118] = 10'b0001000100;
    16'b0000001010000010: out_v[118] = 10'b1110010000;
    16'b0000000010000000: out_v[118] = 10'b1011011011;
    16'b0100000000001000: out_v[118] = 10'b1100101001;
    16'b0100001000000010: out_v[118] = 10'b1000011110;
    16'b0000010000010000: out_v[118] = 10'b1000110100;
    16'b0000011000010000: out_v[118] = 10'b1000011000;
    16'b0000011100010000: out_v[118] = 10'b0010101100;
    16'b0100010100010010: out_v[118] = 10'b0110110100;
    16'b0000010100010010: out_v[118] = 10'b1101000010;
    16'b0000001100010010: out_v[118] = 10'b0101111011;
    16'b0000010100010000: out_v[118] = 10'b0110011000;
    16'b0000000100010010: out_v[118] = 10'b1100110101;
    16'b0100001100010010: out_v[118] = 10'b1001011001;
    16'b0100000100010010: out_v[118] = 10'b0100101000;
    16'b0000001100010000: out_v[118] = 10'b1010011001;
    16'b0000000100010000: out_v[118] = 10'b0010101010;
    16'b0010010000010010: out_v[118] = 10'b0011010001;
    16'b0000010000000011: out_v[118] = 10'b0000100000;
    16'b0110010000000010: out_v[118] = 10'b0000110100;
    16'b0010010000000010: out_v[118] = 10'b1011110000;
    16'b0010010000000000: out_v[118] = 10'b1011111111;
    16'b0000010000000001: out_v[118] = 10'b1011110110;
    16'b0000010100000010: out_v[118] = 10'b0100100101;
    16'b0100010100010000: out_v[118] = 10'b0001111100;
    16'b0000011110010010: out_v[118] = 10'b0111100010;
    16'b0000000000010100: out_v[118] = 10'b0000110011;
    16'b0000000001010100: out_v[118] = 10'b1001011111;
    16'b0000010001010110: out_v[118] = 10'b1111001100;
    16'b0000010101010100: out_v[118] = 10'b0111011111;
    16'b0000000001000100: out_v[118] = 10'b0110110101;
    16'b0000000101010100: out_v[118] = 10'b0111100110;
    16'b0000000100010100: out_v[118] = 10'b0011111111;
    16'b0000000000000100: out_v[118] = 10'b1011011111;
    16'b0000010001010100: out_v[118] = 10'b1001000101;
    16'b0100010000010011: out_v[118] = 10'b0110011010;
    16'b0000010000010011: out_v[118] = 10'b0100100100;
    16'b0100010100000010: out_v[118] = 10'b0111100000;
    16'b0000010001000110: out_v[118] = 10'b1101101001;
    16'b0000000101010110: out_v[118] = 10'b1101010111;
    16'b0000010000010110: out_v[118] = 10'b1111000011;
    16'b0000010101010110: out_v[118] = 10'b1100100111;
    16'b0000000100000010: out_v[118] = 10'b1101101010;
    16'b0000010001000100: out_v[118] = 10'b1001100011;
    default: out_v[118] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000010000000100: out_v[119] = 10'b0111011001;
    16'b0000000010000100: out_v[119] = 10'b1100110011;
    16'b0000010010000101: out_v[119] = 10'b0100100111;
    16'b0010011010000100: out_v[119] = 10'b1011100101;
    16'b0000000010000000: out_v[119] = 10'b1000111001;
    16'b0000010000000000: out_v[119] = 10'b1011000101;
    16'b0000000000000000: out_v[119] = 10'b1101100001;
    16'b0000010010000000: out_v[119] = 10'b1011100101;
    16'b0010001010000000: out_v[119] = 10'b1001010111;
    16'b0000010010000100: out_v[119] = 10'b1110110101;
    16'b0000000000000100: out_v[119] = 10'b0111000111;
    16'b0000001010000100: out_v[119] = 10'b1100101001;
    16'b0010001010000100: out_v[119] = 10'b1001000110;
    16'b0010001010000101: out_v[119] = 10'b0100011101;
    16'b0010011000000100: out_v[119] = 10'b0101000111;
    16'b0010010010000100: out_v[119] = 10'b0100000100;
    16'b0010010000000100: out_v[119] = 10'b1010101011;
    16'b0000001010000101: out_v[119] = 10'b0010001111;
    16'b0100010010000100: out_v[119] = 10'b1111111110;
    16'b0010011000000000: out_v[119] = 10'b0101010111;
    16'b0000011010000100: out_v[119] = 10'b1001110010;
    16'b0100010000000100: out_v[119] = 10'b0101110101;
    16'b0000011000000100: out_v[119] = 10'b1100100010;
    16'b0100000010000000: out_v[119] = 10'b1100110011;
    16'b0010011010000001: out_v[119] = 10'b0000010111;
    16'b0100010000000000: out_v[119] = 10'b0010001001;
    16'b0010000010000100: out_v[119] = 10'b0100010111;
    16'b0010001010000001: out_v[119] = 10'b0010010111;
    16'b0010011010000101: out_v[119] = 10'b0110101001;
    16'b0100000000000000: out_v[119] = 10'b1110101000;
    16'b0010011010000000: out_v[119] = 10'b1000010100;
    16'b0000010110000001: out_v[119] = 10'b0110000111;
    16'b0000010110000000: out_v[119] = 10'b0100100101;
    16'b0000000100000000: out_v[119] = 10'b0000000111;
    16'b0000010100000000: out_v[119] = 10'b1000110011;
    16'b0000000110000000: out_v[119] = 10'b1011100000;
    16'b0010000100000000: out_v[119] = 10'b0111110010;
    16'b0000011110000001: out_v[119] = 10'b0011000100;
    16'b0000000110000001: out_v[119] = 10'b0101010100;
    16'b0000001110000001: out_v[119] = 10'b0101000110;
    16'b0000011110000000: out_v[119] = 10'b1110011100;
    16'b0000000100000001: out_v[119] = 10'b1001001101;
    16'b0000010100000001: out_v[119] = 10'b0110010010;
    16'b0010011110000101: out_v[119] = 10'b1101110111;
    16'b0010000110000000: out_v[119] = 10'b0110111100;
    16'b0000001110000000: out_v[119] = 10'b0011110010;
    16'b0010011110000001: out_v[119] = 10'b0111010110;
    16'b0010001110000001: out_v[119] = 10'b0111000111;
    16'b0010011000000101: out_v[119] = 10'b1001000110;
    16'b0010010010000101: out_v[119] = 10'b0101101011;
    16'b0010000110100001: out_v[119] = 10'b0110000100;
    16'b0010011110000100: out_v[119] = 10'b0000101110;
    16'b0010001110000000: out_v[119] = 10'b1000111000;
    16'b0010010110000001: out_v[119] = 10'b1111000000;
    16'b0010011110000000: out_v[119] = 10'b1010100110;
    16'b0010011000000001: out_v[119] = 10'b1001010110;
    16'b0010000110000001: out_v[119] = 10'b0111010001;
    16'b0000000010000001: out_v[119] = 10'b1000110110;
    16'b0010001110000101: out_v[119] = 10'b1011101100;
    16'b0010001000000001: out_v[119] = 10'b1100010110;
    16'b0010001000000000: out_v[119] = 10'b0111000100;
    16'b0000011010000001: out_v[119] = 10'b0100001010;
    16'b0000000110100001: out_v[119] = 10'b1000111100;
    16'b0010010000000101: out_v[119] = 10'b1010110110;
    16'b0000011010000000: out_v[119] = 10'b1100010000;
    16'b0000011100000000: out_v[119] = 10'b0111011010;
    16'b0000001100000001: out_v[119] = 10'b1111101000;
    16'b0000011110000100: out_v[119] = 10'b0011101000;
    16'b0000011100000100: out_v[119] = 10'b1101100010;
    16'b0010001100000001: out_v[119] = 10'b1011101011;
    16'b0010011100000100: out_v[119] = 10'b0000110111;
    16'b0000001100000000: out_v[119] = 10'b0000111001;
    16'b0010011100000000: out_v[119] = 10'b1100100111;
    16'b0010011100000001: out_v[119] = 10'b1011101000;
    16'b0010000000000000: out_v[119] = 10'b0011101000;
    16'b0000001110000100: out_v[119] = 10'b0001101001;
    16'b0010001100000000: out_v[119] = 10'b1000110011;
    16'b0010001100000100: out_v[119] = 10'b1000010110;
    16'b0000001100000101: out_v[119] = 10'b0011111010;
    16'b0000011100000101: out_v[119] = 10'b0111101010;
    16'b0010010100000000: out_v[119] = 10'b0111001001;
    16'b0010000100000001: out_v[119] = 10'b0011110001;
    16'b0010010100000001: out_v[119] = 10'b0111011001;
    16'b0010010110000000: out_v[119] = 10'b0000101001;
    16'b0000001100000100: out_v[119] = 10'b0110001000;
    16'b0000001000000100: out_v[119] = 10'b0111001110;
    16'b0000011100000001: out_v[119] = 10'b0111111000;
    16'b0010010000000000: out_v[119] = 10'b1101101010;
    16'b0010000000000101: out_v[119] = 10'b1100011111;
    16'b0010001100000101: out_v[119] = 10'b0010011000;
    16'b0010011100000101: out_v[119] = 10'b1100011010;
    16'b0010000100000101: out_v[119] = 10'b1100010101;
    16'b0010001000000101: out_v[119] = 10'b0100010010;
    16'b0010001000000100: out_v[119] = 10'b0011011010;
    16'b0110001000000101: out_v[119] = 10'b1001111011;
    16'b0110001100000101: out_v[119] = 10'b1010010010;
    16'b0010010100000101: out_v[119] = 10'b0000101110;
    16'b0000000000000001: out_v[119] = 10'b1000101010;
    16'b0010010000000001: out_v[119] = 10'b0000100100;
    16'b0000010000000001: out_v[119] = 10'b1010111001;
    16'b0010000000000001: out_v[119] = 10'b1001100001;
    16'b0010000010000001: out_v[119] = 10'b1011101010;
    16'b0010000010000000: out_v[119] = 10'b1011101001;
    16'b0010010010000001: out_v[119] = 10'b1111001010;
    16'b0010010010000000: out_v[119] = 10'b1011011010;
    16'b0000011110000101: out_v[119] = 10'b0001111100;
    16'b0000001110000101: out_v[119] = 10'b0101010010;
    16'b0010001110000100: out_v[119] = 10'b0011001111;
    16'b0000010010000001: out_v[119] = 10'b1111011000;
    16'b0010000010000101: out_v[119] = 10'b0100011110;
    16'b0000001010000000: out_v[119] = 10'b0001001001;
    16'b0000000110000101: out_v[119] = 10'b1011100111;
    16'b0000000110000100: out_v[119] = 10'b1001011000;
    16'b0110001000000100: out_v[119] = 10'b1101100110;
    16'b0010101000000100: out_v[119] = 10'b1111111011;
    16'b0010001000000010: out_v[119] = 10'b0011000111;
    16'b0010101000000000: out_v[119] = 10'b0011000101;
    16'b0010001100000010: out_v[119] = 10'b1100100111;
    16'b0000101000000000: out_v[119] = 10'b0111001101;
    16'b0000001000000000: out_v[119] = 10'b0111001011;
    16'b0010000100000010: out_v[119] = 10'b1101101100;
    16'b0010001000000110: out_v[119] = 10'b0001111110;
    16'b0110001000000110: out_v[119] = 10'b0010111100;
    16'b0000001100000010: out_v[119] = 10'b1010001011;
    16'b0000101100000000: out_v[119] = 10'b1100101011;
    16'b0000000100000010: out_v[119] = 10'b1010000101;
    16'b0010101100000000: out_v[119] = 10'b1001110111;
    16'b0010001100000110: out_v[119] = 10'b1101011111;
    16'b0010001100000011: out_v[119] = 10'b1101000111;
    16'b0010001100000111: out_v[119] = 10'b1101101110;
    16'b0010001000000011: out_v[119] = 10'b1101010011;
    default: out_v[119] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000001010100000: out_v[120] = 10'b1010011011;
    16'b1001000000100100: out_v[120] = 10'b0001011110;
    16'b0000000010100100: out_v[120] = 10'b0110001111;
    16'b0000000000100000: out_v[120] = 10'b0001001001;
    16'b1001000010000000: out_v[120] = 10'b1001001000;
    16'b0101000010100100: out_v[120] = 10'b0100011001;
    16'b1001001010000000: out_v[120] = 10'b0110010011;
    16'b1001000000000100: out_v[120] = 10'b1111010010;
    16'b0000000000100100: out_v[120] = 10'b0010100011;
    16'b1000000010100000: out_v[120] = 10'b1010001111;
    16'b0001000000100000: out_v[120] = 10'b0101100100;
    16'b1101001010100000: out_v[120] = 10'b0010111001;
    16'b0001001000100100: out_v[120] = 10'b1100101001;
    16'b0000000010100000: out_v[120] = 10'b1000001101;
    16'b0100000010100100: out_v[120] = 10'b1010011011;
    16'b1101001000000000: out_v[120] = 10'b0001111110;
    16'b1000001010100000: out_v[120] = 10'b1101010001;
    16'b0001000010100100: out_v[120] = 10'b1001001001;
    16'b0001000000100100: out_v[120] = 10'b1011000011;
    16'b0001000000000100: out_v[120] = 10'b1110110011;
    16'b0000000010000100: out_v[120] = 10'b0101010011;
    16'b0100001010100000: out_v[120] = 10'b0001100110;
    16'b1001000000100000: out_v[120] = 10'b0011100110;
    16'b1101001010000000: out_v[120] = 10'b1011101001;
    16'b1001001010100000: out_v[120] = 10'b1110010001;
    16'b0000000010000000: out_v[120] = 10'b0010011000;
    16'b1001000010100100: out_v[120] = 10'b1001000100;
    16'b0000000000000100: out_v[120] = 10'b1010100001;
    16'b0000001000100000: out_v[120] = 10'b1011111101;
    16'b0101001000100100: out_v[120] = 10'b1101011010;
    16'b0100000000100000: out_v[120] = 10'b0001010101;
    16'b0100001000100100: out_v[120] = 10'b0110011001;
    16'b1001000010100000: out_v[120] = 10'b1000001100;
    16'b0001000000000000: out_v[120] = 10'b1100000101;
    16'b1101001000100100: out_v[120] = 10'b0001011011;
    16'b0100000000100100: out_v[120] = 10'b1001001101;
    16'b0001000010100000: out_v[120] = 10'b0100011000;
    16'b1001001000000000: out_v[120] = 10'b0110110001;
    16'b1001000000000000: out_v[120] = 10'b0111000100;
    16'b0000000000000000: out_v[120] = 10'b0110100011;
    16'b0100000010100000: out_v[120] = 10'b1100100010;
    16'b0000001000100100: out_v[120] = 10'b1001010011;
    16'b1101001000100000: out_v[120] = 10'b1001011010;
    16'b0101000000100100: out_v[120] = 10'b0111100101;
    16'b0100001000100000: out_v[120] = 10'b0101001110;
    16'b1101001010100100: out_v[120] = 10'b0010110011;
    16'b0101000000000000: out_v[120] = 10'b1111100011;
    16'b0101000000100000: out_v[120] = 10'b1011111011;
    16'b0100000000000000: out_v[120] = 10'b0010000110;
    16'b1101000000100000: out_v[120] = 10'b0111100010;
    16'b1101000000000000: out_v[120] = 10'b0110001111;
    16'b0101001000100000: out_v[120] = 10'b0100110001;
    16'b0101001000000000: out_v[120] = 10'b0100011111;
    16'b0100000010000000: out_v[120] = 10'b1010100011;
    16'b1001001000100000: out_v[120] = 10'b0111010101;
    16'b0101000001100000: out_v[120] = 10'b0011010111;
    16'b0101000000100010: out_v[120] = 10'b1101010000;
    16'b1001000010000110: out_v[120] = 10'b0110111011;
    16'b1101000010000000: out_v[120] = 10'b0111000000;
    16'b1001000010000010: out_v[120] = 10'b0111101011;
    16'b1001000000000010: out_v[120] = 10'b0100001101;
    16'b1000000000000100: out_v[120] = 10'b0110010100;
    16'b1001000010000100: out_v[120] = 10'b1000010110;
    16'b1001000010100010: out_v[120] = 10'b0111100110;
    16'b1101000000000110: out_v[120] = 10'b1011110011;
    16'b1100000000000000: out_v[120] = 10'b0100011001;
    16'b1101000000000100: out_v[120] = 10'b1000110011;
    16'b1101000010100000: out_v[120] = 10'b1001011100;
    16'b1100000000000100: out_v[120] = 10'b1100000100;
    16'b1000000010000100: out_v[120] = 10'b0100011010;
    16'b1000000010000000: out_v[120] = 10'b0100010001;
    16'b1101001000000100: out_v[120] = 10'b0000110100;
    16'b1001000011000000: out_v[120] = 10'b1011100111;
    16'b1101000000100100: out_v[120] = 10'b0111110001;
    16'b1000000000000000: out_v[120] = 10'b0100101000;
    16'b1101000000000010: out_v[120] = 10'b1010011010;
    16'b1001000011100000: out_v[120] = 10'b1001001100;
    16'b1001000000100010: out_v[120] = 10'b1010101101;
    16'b1101000000100010: out_v[120] = 10'b1110110010;
    16'b0100000000100010: out_v[120] = 10'b0001110100;
    16'b1100001000100000: out_v[120] = 10'b1100000100;
    16'b0000001000000000: out_v[120] = 10'b0001110011;
    16'b1100001000000000: out_v[120] = 10'b0101010100;
    16'b0100001000000000: out_v[120] = 10'b1000011010;
    16'b1100000000100000: out_v[120] = 10'b1100001001;
    16'b0100001000000100: out_v[120] = 10'b1111011010;
    16'b0100001010100100: out_v[120] = 10'b0101101110;
    16'b1100001010100000: out_v[120] = 10'b0110110001;
    16'b0101001010100100: out_v[120] = 10'b0111111010;
    16'b0101001010100000: out_v[120] = 10'b0001001101;
    16'b1100000010100000: out_v[120] = 10'b1100110001;
    16'b1000000000100000: out_v[120] = 10'b0010111010;
    16'b1000001000100000: out_v[120] = 10'b0000110010;
    16'b0000000011000000: out_v[120] = 10'b1001010011;
    16'b0001001000000000: out_v[120] = 10'b1101010001;
    16'b1000001000000000: out_v[120] = 10'b0111000011;
    16'b0100001010000100: out_v[120] = 10'b1011101100;
    16'b0100001010000000: out_v[120] = 10'b0101100010;
    16'b0001001000100000: out_v[120] = 10'b1111001111;
    16'b1001001000100100: out_v[120] = 10'b0001111010;
    16'b0001001010000000: out_v[120] = 10'b0111010011;
    16'b0001000010100110: out_v[120] = 10'b1111110011;
    16'b1001000000100110: out_v[120] = 10'b1011011111;
    16'b1001000010100110: out_v[120] = 10'b0100001111;
    16'b0001000010000100: out_v[120] = 10'b1001001010;
    16'b0001001000100010: out_v[120] = 10'b1100010111;
    16'b0001000000100110: out_v[120] = 10'b1111011101;
    16'b0101000010100110: out_v[120] = 10'b1111001001;
    16'b0001000010000000: out_v[120] = 10'b0101011000;
    16'b0001001010100000: out_v[120] = 10'b1110100011;
    16'b1001001000100010: out_v[120] = 10'b1101001001;
    16'b0001000000100010: out_v[120] = 10'b1011001100;
    16'b1101000010100110: out_v[120] = 10'b1011101111;
    16'b0001000010100010: out_v[120] = 10'b1011111100;
    16'b1001000000000110: out_v[120] = 10'b1111111111;
    16'b0101000010000000: out_v[120] = 10'b0110111010;
    16'b0101001010000000: out_v[120] = 10'b0100110000;
    16'b1000001010000000: out_v[120] = 10'b1100011000;
    16'b0000001010000000: out_v[120] = 10'b1000010111;
    16'b1100000010000000: out_v[120] = 10'b0110110010;
    default: out_v[120] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000001011010000: out_v[121] = 10'b0110100010;
    16'b0000000010010000: out_v[121] = 10'b1001101011;
    16'b0000101010010001: out_v[121] = 10'b1000110101;
    16'b0000000000010000: out_v[121] = 10'b1100110101;
    16'b0000100000010001: out_v[121] = 10'b1111101100;
    16'b0000100000010000: out_v[121] = 10'b1011000001;
    16'b0000000000000000: out_v[121] = 10'b1000000011;
    16'b0000001000010000: out_v[121] = 10'b1010101010;
    16'b0000100000000000: out_v[121] = 10'b0111011111;
    16'b0000001010010000: out_v[121] = 10'b0010011010;
    16'b0000000011010000: out_v[121] = 10'b0101001101;
    16'b0010000000010000: out_v[121] = 10'b1010110111;
    16'b0000001010010001: out_v[121] = 10'b1000011010;
    16'b0000001010000000: out_v[121] = 10'b0111001001;
    16'b0000101000010001: out_v[121] = 10'b1000000111;
    16'b0010101000010001: out_v[121] = 10'b1000101111;
    16'b0000101010110001: out_v[121] = 10'b1000101110;
    16'b0000001001010000: out_v[121] = 10'b0011010100;
    16'b0000101000010000: out_v[121] = 10'b0011111011;
    16'b0000001011010001: out_v[121] = 10'b0110010001;
    16'b0010101010010001: out_v[121] = 10'b1010100011;
    16'b0010000000000000: out_v[121] = 10'b0100100001;
    16'b0000000001000000: out_v[121] = 10'b0001000110;
    16'b0010001000010000: out_v[121] = 10'b1101010001;
    16'b0000000001010000: out_v[121] = 10'b1101110110;
    16'b0000101010010000: out_v[121] = 10'b0100001101;
    16'b0000101011010001: out_v[121] = 10'b0100110010;
    16'b0010001010010000: out_v[121] = 10'b0010110100;
    16'b0000000010000000: out_v[121] = 10'b0111010101;
    16'b0000001000000000: out_v[121] = 10'b0110000110;
    16'b0000001001000000: out_v[121] = 10'b0011100100;
    16'b0000001001000001: out_v[121] = 10'b0001000110;
    16'b0000001101000000: out_v[121] = 10'b1100101110;
    16'b0000001100010000: out_v[121] = 10'b0000010101;
    16'b0000001111010000: out_v[121] = 10'b1001011111;
    16'b0000001000010001: out_v[121] = 10'b1100001010;
    16'b0000001101010000: out_v[121] = 10'b0000001110;
    16'b0000001011000000: out_v[121] = 10'b1100011000;
    16'b0000001001010001: out_v[121] = 10'b1000011101;
    16'b0000000001000001: out_v[121] = 10'b0011110111;
    16'b0000001110010000: out_v[121] = 10'b0001001000;
    16'b0000001110000000: out_v[121] = 10'b1011001110;
    16'b0000001010000001: out_v[121] = 10'b0111001111;
    16'b0000100001000001: out_v[121] = 10'b1100111001;
    16'b0000100011000001: out_v[121] = 10'b1101001110;
    16'b0000000011000000: out_v[121] = 10'b1100111000;
    16'b0000100010000001: out_v[121] = 10'b1001011010;
    16'b0000100001000101: out_v[121] = 10'b0001111010;
    16'b0000100101000001: out_v[121] = 10'b1001011010;
    16'b0000100000000001: out_v[121] = 10'b0111100000;
    16'b0000000000000001: out_v[121] = 10'b0011011011;
    16'b0010000001010000: out_v[121] = 10'b0100011000;
    16'b0000000010000001: out_v[121] = 10'b1101111100;
    16'b0000101011000001: out_v[121] = 10'b1100100110;
    16'b0000000011000001: out_v[121] = 10'b0110101011;
    16'b0010000001000000: out_v[121] = 10'b0110111010;
    16'b0000101110010001: out_v[121] = 10'b0010110111;
    16'b0000000010010001: out_v[121] = 10'b0000011111;
    16'b0010000010010000: out_v[121] = 10'b0001010011;
    16'b0000101000000001: out_v[121] = 10'b1101110010;
    16'b0000101001000001: out_v[121] = 10'b1001100011;
    16'b0000101001010001: out_v[121] = 10'b1001101011;
    16'b0000100010100001: out_v[121] = 10'b0010010010;
    16'b0000000000010001: out_v[121] = 10'b1011111011;
    16'b0000100010010001: out_v[121] = 10'b0001110001;
    16'b0000000010000011: out_v[121] = 10'b1100000101;
    16'b0000100010110001: out_v[121] = 10'b1001100110;
    16'b0000100000100001: out_v[121] = 10'b0110001001;
    16'b0000000001010001: out_v[121] = 10'b0011100000;
    16'b0000100000110001: out_v[121] = 10'b1111001000;
    16'b0010001011010001: out_v[121] = 10'b1010110110;
    16'b0010001011010000: out_v[121] = 10'b1010111100;
    16'b0010001001010000: out_v[121] = 10'b1100100111;
    16'b0000001011000001: out_v[121] = 10'b0100100011;
    16'b0000101010000001: out_v[121] = 10'b1110100011;
    16'b0000001000000001: out_v[121] = 10'b1001100111;
    16'b0000101001000101: out_v[121] = 10'b1001001010;
    default: out_v[121] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0011010000000000: out_v[122] = 10'b0011001101;
    16'b0011000100000000: out_v[122] = 10'b1100011000;
    16'b0001000100000000: out_v[122] = 10'b0010000111;
    16'b0011010100000000: out_v[122] = 10'b1100011111;
    16'b0011000000000010: out_v[122] = 10'b0010011101;
    16'b0001000000000000: out_v[122] = 10'b0000100001;
    16'b0000000100000000: out_v[122] = 10'b1011110011;
    16'b0010010000000010: out_v[122] = 10'b1000100111;
    16'b0000000000000000: out_v[122] = 10'b0111001100;
    16'b1011010000000010: out_v[122] = 10'b0000011011;
    16'b1001000000000000: out_v[122] = 10'b0100110001;
    16'b0011000000000000: out_v[122] = 10'b1000000111;
    16'b0011010000000010: out_v[122] = 10'b0010110111;
    16'b1001000100000000: out_v[122] = 10'b1001100011;
    16'b1000000000000000: out_v[122] = 10'b0000001110;
    16'b0001000000000010: out_v[122] = 10'b1111100110;
    16'b1011000000000000: out_v[122] = 10'b0111001011;
    16'b0010010000000000: out_v[122] = 10'b1100100011;
    16'b0010010100000000: out_v[122] = 10'b0000110001;
    16'b1011000100000000: out_v[122] = 10'b1001010111;
    16'b0011000100000010: out_v[122] = 10'b0101001000;
    16'b0011010100000010: out_v[122] = 10'b0110100001;
    16'b1011010000000000: out_v[122] = 10'b0101101000;
    16'b1011010100000000: out_v[122] = 10'b1100011011;
    16'b1011000000000010: out_v[122] = 10'b0110010111;
    16'b0000010000000000: out_v[122] = 10'b0100101101;
    16'b1000010000000000: out_v[122] = 10'b1000111010;
    16'b1000000000000010: out_v[122] = 10'b0111110010;
    16'b1000010000000010: out_v[122] = 10'b1000001011;
    16'b1001010000000000: out_v[122] = 10'b0100011110;
    16'b1000001000000000: out_v[122] = 10'b0000001001;
    16'b0000000000000010: out_v[122] = 10'b0011111000;
    16'b0000011000000010: out_v[122] = 10'b1100010110;
    16'b0000010000000010: out_v[122] = 10'b0010010001;
    16'b1000000100000000: out_v[122] = 10'b0110001110;
    16'b1000011000000000: out_v[122] = 10'b1011001011;
    16'b0000011000000000: out_v[122] = 10'b0010111110;
    16'b0010011000000010: out_v[122] = 10'b0010100110;
    16'b0000010100000010: out_v[122] = 10'b0010001110;
    16'b0001000100000010: out_v[122] = 10'b1111001100;
    16'b0010010100000010: out_v[122] = 10'b0111110110;
    16'b0011011000000010: out_v[122] = 10'b0001010100;
    16'b0000001000000010: out_v[122] = 10'b0001000110;
    16'b0011011000000000: out_v[122] = 10'b1111011011;
    16'b1000001000000010: out_v[122] = 10'b0011001001;
    16'b1000010100000000: out_v[122] = 10'b1010100010;
    16'b1000000100000010: out_v[122] = 10'b1100111111;
    16'b0000010100000000: out_v[122] = 10'b0110001011;
    16'b0000000100000010: out_v[122] = 10'b0001100110;
    16'b1011011000000000: out_v[122] = 10'b1001111110;
    16'b1010010000000000: out_v[122] = 10'b1001101010;
    16'b1011010100000010: out_v[122] = 10'b1000011100;
    16'b1010011000000000: out_v[122] = 10'b1010111010;
    16'b1010010100000000: out_v[122] = 10'b0101110000;
    16'b1001010000000010: out_v[122] = 10'b1100001010;
    16'b1000010100000010: out_v[122] = 10'b1000111110;
    16'b1010010000000010: out_v[122] = 10'b1100000100;
    16'b0011110100000010: out_v[122] = 10'b1111010010;
    16'b0000110100000010: out_v[122] = 10'b0111101110;
    16'b0000100000000010: out_v[122] = 10'b0101010011;
    16'b0000110000000010: out_v[122] = 10'b0111010011;
    16'b0011110000000010: out_v[122] = 10'b0011110111;
    16'b1001000000000010: out_v[122] = 10'b1000110100;
    16'b0000100100000000: out_v[122] = 10'b0100101010;
    16'b0000100100000010: out_v[122] = 10'b0111101110;
    16'b0011011100000010: out_v[122] = 10'b1100001111;
    16'b0000001100000010: out_v[122] = 10'b1011100111;
    16'b1011110100000010: out_v[122] = 10'b1100011100;
    16'b0011110100000000: out_v[122] = 10'b0110011110;
    16'b0010110100000010: out_v[122] = 10'b0110001011;
    16'b0011010100001010: out_v[122] = 10'b1010000111;
    16'b0010110100000000: out_v[122] = 10'b0011011111;
    16'b1000100100000010: out_v[122] = 10'b1011101001;
    16'b1001010100000010: out_v[122] = 10'b1111001011;
    16'b1010010100000010: out_v[122] = 10'b1011100111;
    16'b1000110100000010: out_v[122] = 10'b1001100111;
    16'b1000110000000010: out_v[122] = 10'b0101110100;
    16'b1000100000000010: out_v[122] = 10'b1011001001;
    16'b1010110100000010: out_v[122] = 10'b1110000011;
    16'b0011010101000010: out_v[122] = 10'b0001101111;
    16'b0010010101000010: out_v[122] = 10'b0111001011;
    16'b0000010101000010: out_v[122] = 10'b0011111110;
    16'b0010110000000010: out_v[122] = 10'b1000110110;
    default: out_v[122] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1000000100000100: out_v[123] = 10'b1111000101;
    16'b1000100110100000: out_v[123] = 10'b1011000011;
    16'b1000100010100000: out_v[123] = 10'b0010110011;
    16'b0000000010000000: out_v[123] = 10'b0110010111;
    16'b0000000110000000: out_v[123] = 10'b0100101101;
    16'b1000000100000001: out_v[123] = 10'b1111000001;
    16'b1000000000000000: out_v[123] = 10'b0010001010;
    16'b1000100010000000: out_v[123] = 10'b1100110111;
    16'b1000000010000000: out_v[123] = 10'b0100110101;
    16'b0000100010000000: out_v[123] = 10'b1100110101;
    16'b1000100110000000: out_v[123] = 10'b0101011001;
    16'b1000000010000001: out_v[123] = 10'b0010110111;
    16'b1000100000000000: out_v[123] = 10'b1010101001;
    16'b1000100010100100: out_v[123] = 10'b1101000011;
    16'b0000000000000100: out_v[123] = 10'b0011110100;
    16'b0000000000000000: out_v[123] = 10'b0001110011;
    16'b1000000110000000: out_v[123] = 10'b0010111011;
    16'b1000100010000001: out_v[123] = 10'b0010101110;
    16'b1000000110000001: out_v[123] = 10'b1101100010;
    16'b1000000010000100: out_v[123] = 10'b1111111110;
    16'b1000000100000000: out_v[123] = 10'b0101000100;
    16'b0000000010000100: out_v[123] = 10'b0110011011;
    16'b0000100010100100: out_v[123] = 10'b1101100101;
    16'b1000100010000100: out_v[123] = 10'b0110010110;
    16'b0000000000000001: out_v[123] = 10'b0010010011;
    16'b0000000010100100: out_v[123] = 10'b1000110111;
    16'b1000000010100100: out_v[123] = 10'b1111010010;
    16'b1000000000000001: out_v[123] = 10'b1000011000;
    16'b0000000100000001: out_v[123] = 10'b1001001110;
    16'b0000000100000000: out_v[123] = 10'b0001000101;
    16'b1000000110000100: out_v[123] = 10'b1101010111;
    16'b0000100010000100: out_v[123] = 10'b1011001011;
    16'b0000000010000001: out_v[123] = 10'b0101001010;
    16'b1000100110000001: out_v[123] = 10'b0100001111;
    16'b0000110100000001: out_v[123] = 10'b1110100011;
    16'b0000010000000001: out_v[123] = 10'b0100110110;
    16'b0000010000000100: out_v[123] = 10'b0111011000;
    16'b1000010000000100: out_v[123] = 10'b0111000111;
    16'b1000010000000000: out_v[123] = 10'b1111000011;
    16'b0000010000000000: out_v[123] = 10'b1101000011;
    16'b0000110100100001: out_v[123] = 10'b1111010111;
    16'b0000010100000001: out_v[123] = 10'b0000101100;
    16'b0000110000000001: out_v[123] = 10'b0110010000;
    16'b1000010100000000: out_v[123] = 10'b1111011010;
    16'b1000010000000101: out_v[123] = 10'b0111000110;
    16'b0000010100000000: out_v[123] = 10'b1110110100;
    16'b1000010000000001: out_v[123] = 10'b0111010101;
    16'b1000010100000001: out_v[123] = 10'b0001100110;
    16'b1000010100000100: out_v[123] = 10'b1010011010;
    16'b0000010000100001: out_v[123] = 10'b0010110110;
    16'b0000110110100001: out_v[123] = 10'b0000101010;
    16'b0000110110000001: out_v[123] = 10'b0000011111;
    16'b0000110000100001: out_v[123] = 10'b1001000111;
    16'b1000000000000100: out_v[123] = 10'b1000001010;
    16'b1000010100000101: out_v[123] = 10'b0010110011;
    16'b0000110010000000: out_v[123] = 10'b0111101100;
    16'b0000010000000101: out_v[123] = 10'b0101010101;
    16'b0010010100000001: out_v[123] = 10'b0001001111;
    16'b0010000000000001: out_v[123] = 10'b1001001100;
    16'b0000010010000001: out_v[123] = 10'b1100100110;
    16'b0000110010000001: out_v[123] = 10'b1000100111;
    16'b0000010110000000: out_v[123] = 10'b0010100110;
    16'b0000100110000000: out_v[123] = 10'b0001010111;
    16'b0000110110000000: out_v[123] = 10'b0011010110;
    16'b0000010110000001: out_v[123] = 10'b0001111011;
    16'b0000100010000001: out_v[123] = 10'b0100011011;
    16'b0000100110000001: out_v[123] = 10'b1100011101;
    16'b0010010000000001: out_v[123] = 10'b1001010110;
    16'b1010010100000000: out_v[123] = 10'b0010110111;
    16'b0010010100000000: out_v[123] = 10'b1110011110;
    16'b1000110110000001: out_v[123] = 10'b0110011110;
    16'b1000110110000000: out_v[123] = 10'b0011110110;
    16'b0000000000100101: out_v[123] = 10'b0001100101;
    16'b1000000000100100: out_v[123] = 10'b1011010110;
    16'b0000000000000101: out_v[123] = 10'b1011010001;
    16'b0000000100100101: out_v[123] = 10'b0110110111;
    16'b0000010100000101: out_v[123] = 10'b1101001010;
    16'b0000000100000101: out_v[123] = 10'b1011100010;
    16'b1000000000000101: out_v[123] = 10'b1000100010;
    16'b1000000000100001: out_v[123] = 10'b1011101100;
    16'b0000010100000100: out_v[123] = 10'b0100111010;
    16'b0000000100000100: out_v[123] = 10'b0101110101;
    16'b1000000100000101: out_v[123] = 10'b1111000101;
    16'b0000010100100101: out_v[123] = 10'b0001011001;
    16'b1000000100100101: out_v[123] = 10'b0010001011;
    16'b1010000000000001: out_v[123] = 10'b0011011010;
    16'b0000100000000001: out_v[123] = 10'b0000111010;
    16'b1000100000000001: out_v[123] = 10'b0111100110;
    16'b1010000000000000: out_v[123] = 10'b0001001000;
    16'b0000010100100001: out_v[123] = 10'b0011101001;
    16'b0010000100000001: out_v[123] = 10'b1001111111;
    16'b0000000100100001: out_v[123] = 10'b0000010111;
    16'b1000000000100101: out_v[123] = 10'b0101011010;
    16'b0000000000100001: out_v[123] = 10'b1101010011;
    16'b0000110110100101: out_v[123] = 10'b0100001101;
    16'b0000100110100001: out_v[123] = 10'b0011001110;
    16'b1010000100000001: out_v[123] = 10'b1110100010;
    16'b0000110100000101: out_v[123] = 10'b0011011001;
    16'b0000100110000101: out_v[123] = 10'b1101011110;
    16'b1000110100000101: out_v[123] = 10'b1111000101;
    16'b0000010110000101: out_v[123] = 10'b1110111011;
    16'b1000010110000001: out_v[123] = 10'b0110011001;
    16'b1000110100000001: out_v[123] = 10'b0100110000;
    16'b1000010110000000: out_v[123] = 10'b1001110100;
    16'b0000000110000101: out_v[123] = 10'b1100000100;
    16'b0000110110000101: out_v[123] = 10'b0110001111;
    16'b1000110110100001: out_v[123] = 10'b1100010010;
    16'b1000110110000101: out_v[123] = 10'b0101011100;
    16'b0000110110000100: out_v[123] = 10'b1000010010;
    16'b0000100000000101: out_v[123] = 10'b0011110011;
    16'b1000010110000100: out_v[123] = 10'b0011111111;
    16'b0000100100000100: out_v[123] = 10'b0111101110;
    16'b1000110100000100: out_v[123] = 10'b1010100101;
    16'b0000100000100101: out_v[123] = 10'b1010010111;
    16'b1000110100100000: out_v[123] = 10'b0011110001;
    16'b1000110110100000: out_v[123] = 10'b1000101110;
    16'b1000110100000000: out_v[123] = 10'b0001101010;
    16'b1000110100100100: out_v[123] = 10'b1010010111;
    16'b1000100100000000: out_v[123] = 10'b0111011101;
    16'b1000100000100101: out_v[123] = 10'b1110111010;
    16'b0000110100100100: out_v[123] = 10'b1111100110;
    16'b0000110100000000: out_v[123] = 10'b1111111000;
    16'b0000100100100100: out_v[123] = 10'b1011110101;
    16'b1000110110000100: out_v[123] = 10'b1011111011;
    16'b1000110110100100: out_v[123] = 10'b1010111010;
    16'b0000100100000101: out_v[123] = 10'b0011111010;
    16'b0000100000000100: out_v[123] = 10'b0111111111;
    16'b0000100100000000: out_v[123] = 10'b1011010110;
    16'b1000100100100100: out_v[123] = 10'b1001001011;
    16'b0000100000000000: out_v[123] = 10'b1001100101;
    16'b0000100100000001: out_v[123] = 10'b0100100110;
    16'b1000100100000100: out_v[123] = 10'b1110110111;
    16'b0000110100000100: out_v[123] = 10'b1010101110;
    16'b1000100100000001: out_v[123] = 10'b0011110100;
    16'b1000100000000101: out_v[123] = 10'b1011100100;
    16'b0000100000100100: out_v[123] = 10'b1011111010;
    16'b1000010110100000: out_v[123] = 10'b1001100011;
    16'b1000100100100000: out_v[123] = 10'b1110001110;
    16'b1000000010100001: out_v[123] = 10'b1101100101;
    16'b1000000010000101: out_v[123] = 10'b0000101000;
    16'b1000000010100000: out_v[123] = 10'b0010111110;
    16'b1000110010100001: out_v[123] = 10'b0011011001;
    16'b0000000010100001: out_v[123] = 10'b1110100110;
    16'b0000000010000101: out_v[123] = 10'b1010001101;
    16'b1000010010000001: out_v[123] = 10'b1111000011;
    16'b0000010010100001: out_v[123] = 10'b1001010111;
    16'b1000010010100001: out_v[123] = 10'b0010010001;
    16'b0000000010100000: out_v[123] = 10'b0011101001;
    16'b1000010010000101: out_v[123] = 10'b0011110010;
    16'b1000010110000101: out_v[123] = 10'b0101011000;
    16'b1000110110100101: out_v[123] = 10'b0010011110;
    16'b0000010110100101: out_v[123] = 10'b0101101101;
    16'b1000010110100001: out_v[123] = 10'b1101010101;
    16'b0000010010000101: out_v[123] = 10'b1110000111;
    16'b1000010110100101: out_v[123] = 10'b1101011010;
    16'b0000000110000001: out_v[123] = 10'b0100010110;
    16'b1000000110100001: out_v[123] = 10'b0111100011;
    16'b1000000110000101: out_v[123] = 10'b0111010101;
    default: out_v[123] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1100100001000010: out_v[124] = 10'b1101000010;
    16'b1000100011001010: out_v[124] = 10'b0010111001;
    16'b1101000000001110: out_v[124] = 10'b1101101100;
    16'b1100100001001010: out_v[124] = 10'b0111101110;
    16'b1101000000001100: out_v[124] = 10'b1100111101;
    16'b1100000011001011: out_v[124] = 10'b0100100110;
    16'b1101000000001000: out_v[124] = 10'b0100001001;
    16'b1000100001001010: out_v[124] = 10'b1010011001;
    16'b1100000000001010: out_v[124] = 10'b1110111101;
    16'b1100100011001010: out_v[124] = 10'b0110100010;
    16'b1100000011001010: out_v[124] = 10'b0010100001;
    16'b1100100001001110: out_v[124] = 10'b1110001010;
    16'b1100000001001010: out_v[124] = 10'b1000101001;
    16'b1100000001001110: out_v[124] = 10'b0111001010;
    16'b0100000001001010: out_v[124] = 10'b0110010101;
    16'b1100000000001000: out_v[124] = 10'b0011010111;
    16'b0101000000100100: out_v[124] = 10'b1111110010;
    16'b0101000000000000: out_v[124] = 10'b1110100110;
    16'b1101000001001110: out_v[124] = 10'b0111110111;
    16'b0000100001001010: out_v[124] = 10'b1011000111;
    16'b1100000010001010: out_v[124] = 10'b1101101101;
    16'b0001000000000100: out_v[124] = 10'b1011011011;
    16'b1101000010001100: out_v[124] = 10'b1111111110;
    16'b1100000000000000: out_v[124] = 10'b1010101001;
    16'b1101000001001010: out_v[124] = 10'b0111111000;
    16'b0100000011001010: out_v[124] = 10'b0011100001;
    16'b1101000010001010: out_v[124] = 10'b0001110110;
    16'b1101000000001010: out_v[124] = 10'b1101110111;
    16'b1100000001000010: out_v[124] = 10'b0010100101;
    16'b0000100000001000: out_v[124] = 10'b0111100011;
    16'b0100100001001010: out_v[124] = 10'b0001011111;
    16'b1101000010001110: out_v[124] = 10'b0111000011;
    16'b1111000000001100: out_v[124] = 10'b1011100111;
    16'b1101000000000100: out_v[124] = 10'b1010101110;
    16'b1100100001001011: out_v[124] = 10'b0000001011;
    16'b0101000000000100: out_v[124] = 10'b1011100100;
    16'b0101000000001100: out_v[124] = 10'b1000010111;
    16'b1100100000001010: out_v[124] = 10'b0111011110;
    16'b1110100001001010: out_v[124] = 10'b1110110110;
    16'b0000100000000001: out_v[124] = 10'b1010100010;
    16'b0000000000000001: out_v[124] = 10'b1001100111;
    16'b0000000000001000: out_v[124] = 10'b0010111000;
    16'b0000000000000000: out_v[124] = 10'b0110111000;
    16'b0000000000001001: out_v[124] = 10'b0100001001;
    16'b0000000010000001: out_v[124] = 10'b0001111011;
    16'b0010000000001000: out_v[124] = 10'b0011001011;
    16'b0100000000001000: out_v[124] = 10'b1001110110;
    16'b0000100010000001: out_v[124] = 10'b0011001011;
    16'b0000100000001001: out_v[124] = 10'b1001001100;
    16'b0010000000001001: out_v[124] = 10'b1000100101;
    16'b1010000000001001: out_v[124] = 10'b1010100100;
    16'b1000100000000011: out_v[124] = 10'b0001111000;
    16'b1000100000000001: out_v[124] = 10'b1101001001;
    16'b0010100000101001: out_v[124] = 10'b0110110111;
    16'b1010100001001011: out_v[124] = 10'b1100111110;
    16'b1010100001001010: out_v[124] = 10'b0000110110;
    16'b0001100001000011: out_v[124] = 10'b1011100110;
    16'b0010100000000001: out_v[124] = 10'b1000101111;
    16'b0010100000001001: out_v[124] = 10'b0000111011;
    16'b1010100000001000: out_v[124] = 10'b1001010100;
    16'b1010100000101001: out_v[124] = 10'b1101010110;
    16'b1000100001000011: out_v[124] = 10'b0011010011;
    16'b1010100000001001: out_v[124] = 10'b1010100011;
    16'b0010000000000001: out_v[124] = 10'b0001100100;
    16'b0010000000001101: out_v[124] = 10'b1110111101;
    16'b1000100000001001: out_v[124] = 10'b0010110101;
    16'b0100000000001101: out_v[124] = 10'b0101010011;
    16'b0100000000001001: out_v[124] = 10'b0100100101;
    16'b1010100001101011: out_v[124] = 10'b1101011011;
    16'b0010100000001000: out_v[124] = 10'b1010000100;
    16'b0000100010001001: out_v[124] = 10'b1011100100;
    16'b1000100001001011: out_v[124] = 10'b1100001011;
    16'b1010100000000001: out_v[124] = 10'b1111111100;
    16'b0010100000101000: out_v[124] = 10'b1101110111;
    16'b0000000000001101: out_v[124] = 10'b1001011011;
    16'b0100100000001001: out_v[124] = 10'b1000101100;
    16'b1000100011000011: out_v[124] = 10'b1001100111;
    16'b1000000001000110: out_v[124] = 10'b1001110010;
    16'b1010000000001010: out_v[124] = 10'b0011111001;
    16'b0000000001001010: out_v[124] = 10'b0110101101;
    16'b1000000001000010: out_v[124] = 10'b0011011001;
    16'b1010000001001010: out_v[124] = 10'b1110110010;
    16'b1000000000000010: out_v[124] = 10'b0110111001;
    16'b1000100001000010: out_v[124] = 10'b1101010011;
    16'b1000000011001010: out_v[124] = 10'b0110001101;
    16'b1000000001001010: out_v[124] = 10'b0010110100;
    16'b1000000000000000: out_v[124] = 10'b0110011101;
    16'b1000000000000110: out_v[124] = 10'b1001101011;
    16'b1110000001001010: out_v[124] = 10'b0011011001;
    16'b1000100001001110: out_v[124] = 10'b1000101010;
    16'b0000000000001010: out_v[124] = 10'b0011111110;
    16'b1000000000001010: out_v[124] = 10'b0101000101;
    16'b1000100000000010: out_v[124] = 10'b0111101110;
    16'b1010000001000010: out_v[124] = 10'b1011111100;
    16'b1000000000001000: out_v[124] = 10'b1000010111;
    16'b1010000000000000: out_v[124] = 10'b1001001011;
    16'b0000000010001000: out_v[124] = 10'b1010110010;
    16'b1000100000001010: out_v[124] = 10'b1001011001;
    16'b1000100001000110: out_v[124] = 10'b1011000000;
    16'b1000000001001110: out_v[124] = 10'b1111001100;
    16'b1010000000001000: out_v[124] = 10'b1101001001;
    16'b1100000001000110: out_v[124] = 10'b0011010100;
    16'b0000000001000010: out_v[124] = 10'b0011001010;
    16'b1010000000000010: out_v[124] = 10'b1011001111;
    16'b0100100001001111: out_v[124] = 10'b1000110110;
    16'b0100000000000000: out_v[124] = 10'b1001010110;
    16'b0100100001001000: out_v[124] = 10'b0001001011;
    16'b0100100011001010: out_v[124] = 10'b1100100100;
    16'b1000100001000111: out_v[124] = 10'b1000011001;
    16'b0100100001000011: out_v[124] = 10'b0111111110;
    16'b0000000000001100: out_v[124] = 10'b1000010010;
    16'b0100100000000001: out_v[124] = 10'b1101111000;
    16'b0100100000000000: out_v[124] = 10'b1100000001;
    16'b0100100000001000: out_v[124] = 10'b1110000011;
    16'b0100000000001100: out_v[124] = 10'b1011110110;
    16'b0100100010001000: out_v[124] = 10'b1110100101;
    16'b0000100000000100: out_v[124] = 10'b1011011111;
    16'b0100100011001011: out_v[124] = 10'b1011100111;
    16'b1100100001000110: out_v[124] = 10'b1001100111;
    16'b0100100010000001: out_v[124] = 10'b1001111110;
    16'b0000100000000000: out_v[124] = 10'b1100100111;
    16'b0100000010000001: out_v[124] = 10'b0111011000;
    16'b0100100011000011: out_v[124] = 10'b0110011100;
    16'b0000100001000011: out_v[124] = 10'b0001100111;
    16'b0000100001001110: out_v[124] = 10'b0100010111;
    16'b0100100011001000: out_v[124] = 10'b0010010111;
    16'b0100100001001011: out_v[124] = 10'b0001111010;
    16'b1100100001000111: out_v[124] = 10'b1001101010;
    16'b0100000000000001: out_v[124] = 10'b1011000101;
    16'b0100100001001110: out_v[124] = 10'b0011100111;
    16'b0100100001000010: out_v[124] = 10'b1101010110;
    16'b0100100000001100: out_v[124] = 10'b0011110111;
    16'b1100100001000011: out_v[124] = 10'b1000010001;
    16'b0101100001001010: out_v[124] = 10'b1001111111;
    16'b0000100000001100: out_v[124] = 10'b1100000101;
    16'b0100100011001110: out_v[124] = 10'b0100101010;
    16'b1100000011000110: out_v[124] = 10'b1011101111;
    16'b1100000011001110: out_v[124] = 10'b1000011111;
    16'b0100000010001000: out_v[124] = 10'b0001111111;
    16'b1100000011000010: out_v[124] = 10'b0001100111;
    16'b0100100010001001: out_v[124] = 10'b1100101001;
    16'b0000100010001000: out_v[124] = 10'b1111100100;
    16'b1100000000000010: out_v[124] = 10'b1111110110;
    16'b0000000010001001: out_v[124] = 10'b1000110100;
    16'b1111100001001111: out_v[124] = 10'b0000110111;
    16'b1111100001001011: out_v[124] = 10'b1101100110;
    16'b1101100000001011: out_v[124] = 10'b1011011100;
    16'b1000100000001011: out_v[124] = 10'b1011110010;
    16'b1110100001001011: out_v[124] = 10'b0011001011;
    16'b1101100000001001: out_v[124] = 10'b0011101011;
    16'b1100100000001011: out_v[124] = 10'b0001111101;
    16'b0000100001001011: out_v[124] = 10'b1011111010;
    16'b1100100000001001: out_v[124] = 10'b0100011001;
    16'b1100000001001011: out_v[124] = 10'b0111000010;
    16'b1101100001001011: out_v[124] = 10'b0111010010;
    16'b1111100000001101: out_v[124] = 10'b1011011010;
    16'b1111100000001001: out_v[124] = 10'b1110011110;
    16'b1110100001001111: out_v[124] = 10'b0011010111;
    16'b0100000001001110: out_v[124] = 10'b1100100111;
    16'b0100000001001111: out_v[124] = 10'b1010001100;
    16'b0100000000000101: out_v[124] = 10'b1011000110;
    16'b0100000001001100: out_v[124] = 10'b1010110010;
    16'b0100000000000100: out_v[124] = 10'b0011111101;
    16'b0100000001001000: out_v[124] = 10'b1001011011;
    16'b0000000001001110: out_v[124] = 10'b1111011011;
    16'b0100000001001101: out_v[124] = 10'b0111110101;
    16'b0100000010001001: out_v[124] = 10'b0101100100;
    16'b1100000000000001: out_v[124] = 10'b0110010001;
    16'b0100100000001101: out_v[124] = 10'b0100110000;
    16'b1100000000000101: out_v[124] = 10'b0100011001;
    16'b1100000000000111: out_v[124] = 10'b0110010111;
    16'b1100100001001111: out_v[124] = 10'b1011001001;
    16'b0100100010001101: out_v[124] = 10'b1100001001;
    16'b0100100000000101: out_v[124] = 10'b0011011110;
    16'b0100100001001001: out_v[124] = 10'b1001011111;
    default: out_v[124] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1100010000010001: out_v[125] = 10'b0111000011;
    16'b0100110000000001: out_v[125] = 10'b0100100101;
    16'b1100110000001001: out_v[125] = 10'b1110011100;
    16'b0100100000001001: out_v[125] = 10'b1001010101;
    16'b1000000000010001: out_v[125] = 10'b0010100101;
    16'b1000110000000001: out_v[125] = 10'b0010110011;
    16'b1000111000001001: out_v[125] = 10'b0111101100;
    16'b1000110000001001: out_v[125] = 10'b0101000111;
    16'b0100101000001001: out_v[125] = 10'b1101011011;
    16'b1100000000000001: out_v[125] = 10'b1011110010;
    16'b1000111000001000: out_v[125] = 10'b1100010011;
    16'b1100110000000001: out_v[125] = 10'b0011110001;
    16'b0100100000000001: out_v[125] = 10'b0111001101;
    16'b0100000000000001: out_v[125] = 10'b1000101000;
    16'b0000100000001001: out_v[125] = 10'b1001101011;
    16'b1000110000000000: out_v[125] = 10'b0101001000;
    16'b1100100000001001: out_v[125] = 10'b0010111111;
    16'b0000000000000001: out_v[125] = 10'b0100011011;
    16'b1000111000011000: out_v[125] = 10'b0001111001;
    16'b1000101000001001: out_v[125] = 10'b1101100111;
    16'b0000101000001001: out_v[125] = 10'b0111111010;
    16'b0100111000001001: out_v[125] = 10'b1111010111;
    16'b1000100000001001: out_v[125] = 10'b0011101111;
    16'b0000100000000001: out_v[125] = 10'b1101000110;
    16'b0100110000001001: out_v[125] = 10'b1000111011;
    16'b1000100000000001: out_v[125] = 10'b1000111111;
    16'b1000110000011000: out_v[125] = 10'b1101001011;
    16'b0100010000000001: out_v[125] = 10'b1000101010;
    16'b0000110000000001: out_v[125] = 10'b0101000001;
    16'b1000110000001000: out_v[125] = 10'b1000111111;
    16'b1100100000000001: out_v[125] = 10'b0010111011;
    16'b1100101000001001: out_v[125] = 10'b0111100110;
    16'b0100000000001001: out_v[125] = 10'b0010010110;
    16'b1000000000000001: out_v[125] = 10'b0001101100;
    16'b1000000000010000: out_v[125] = 10'b0111011000;
    16'b1100010000000001: out_v[125] = 10'b0010011100;
    16'b0000110000001001: out_v[125] = 10'b1001111111;
    16'b1100111000001001: out_v[125] = 10'b1111110101;
    16'b1000110000010000: out_v[125] = 10'b1011110100;
    16'b1000110000010001: out_v[125] = 10'b0011011110;
    16'b1000101000001000: out_v[125] = 10'b0011111000;
    16'b1100110000010001: out_v[125] = 10'b0001110011;
    16'b0100101000000001: out_v[125] = 10'b1100010110;
    16'b1000010000010001: out_v[125] = 10'b1101100100;
    16'b1100000000010001: out_v[125] = 10'b0110000011;
    16'b0000010000000000: out_v[125] = 10'b1101000100;
    16'b1000010000000000: out_v[125] = 10'b0100101010;
    16'b1000010000010000: out_v[125] = 10'b0111000001;
    16'b1000010000000001: out_v[125] = 10'b1110101000;
    16'b1000000000000000: out_v[125] = 10'b0111001011;
    16'b0000010000000001: out_v[125] = 10'b1000111010;
    16'b0000000000000000: out_v[125] = 10'b0100110111;
    16'b1000010000010011: out_v[125] = 10'b0110011100;
    16'b1000100000000011: out_v[125] = 10'b1111110010;
    16'b1000010000010010: out_v[125] = 10'b1101000101;
    16'b1100000000010011: out_v[125] = 10'b1101110110;
    16'b1000100000010001: out_v[125] = 10'b1010011001;
    16'b1000100000000000: out_v[125] = 10'b1001110110;
    16'b1000000000010011: out_v[125] = 10'b1111010100;
    16'b1000010000110000: out_v[125] = 10'b1000010111;
    16'b0100000000000011: out_v[125] = 10'b0010101011;
    16'b1000100000110000: out_v[125] = 10'b1011111111;
    16'b1000100000000010: out_v[125] = 10'b1100010110;
    16'b1000000000010010: out_v[125] = 10'b1011000101;
    16'b1000100000010000: out_v[125] = 10'b1000110100;
    16'b0000100000000011: out_v[125] = 10'b0100000100;
    16'b1000100000010010: out_v[125] = 10'b0011011010;
    16'b1100000000000011: out_v[125] = 10'b1111110101;
    16'b0000100000000000: out_v[125] = 10'b0010000011;
    16'b1000000000110000: out_v[125] = 10'b0001011111;
    16'b1000000000000011: out_v[125] = 10'b1110110000;
    16'b0000000000000011: out_v[125] = 10'b1001100010;
    16'b1000011000010000: out_v[125] = 10'b0000111101;
    16'b0100010000000011: out_v[125] = 10'b1000001111;
    16'b0100000000000000: out_v[125] = 10'b0000100101;
    16'b0100010000000000: out_v[125] = 10'b1011000000;
    16'b1000010000000011: out_v[125] = 10'b1011011010;
    16'b1100010000000011: out_v[125] = 10'b1111011010;
    16'b1000010000000010: out_v[125] = 10'b1000110100;
    16'b0000010000000011: out_v[125] = 10'b0000011010;
    16'b0000100000001000: out_v[125] = 10'b0000110001;
    16'b1000100000011000: out_v[125] = 10'b1001110000;
    16'b0000000000001000: out_v[125] = 10'b0010011000;
    16'b0000110000001000: out_v[125] = 10'b1010011010;
    16'b0000101000001000: out_v[125] = 10'b0101110010;
    16'b0000000000010000: out_v[125] = 10'b1010111010;
    16'b0000110000000000: out_v[125] = 10'b0110000000;
    16'b0001100000001000: out_v[125] = 10'b1001110000;
    16'b0000100000011000: out_v[125] = 10'b1000100110;
    16'b0000100000010000: out_v[125] = 10'b1010110011;
    16'b0000110000010000: out_v[125] = 10'b1100110011;
    16'b0100010000001001: out_v[125] = 10'b1001100010;
    16'b1000101000011010: out_v[125] = 10'b0011000011;
    16'b1000101000000000: out_v[125] = 10'b1101010110;
    16'b1000101000011000: out_v[125] = 10'b0111101001;
    16'b1000100000011010: out_v[125] = 10'b0000110010;
    16'b1000100000001000: out_v[125] = 10'b1011001011;
    16'b1000101000010000: out_v[125] = 10'b1100001111;
    16'b0001010000000000: out_v[125] = 10'b0111110010;
    16'b0001000000000000: out_v[125] = 10'b0010101011;
    16'b0000010000001000: out_v[125] = 10'b1111001101;
    16'b0001010000001000: out_v[125] = 10'b0110000100;
    16'b1100010000001001: out_v[125] = 10'b0101011110;
    16'b0101010000000001: out_v[125] = 10'b0001110111;
    16'b1100000000010000: out_v[125] = 10'b0110010001;
    16'b0100000000010001: out_v[125] = 10'b1000001000;
    16'b1100010000010000: out_v[125] = 10'b0000101000;
    default: out_v[125] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000000010000: out_v[126] = 10'b1010100010;
    16'b0100000000010000: out_v[126] = 10'b1111001110;
    16'b0100000000010110: out_v[126] = 10'b0010000111;
    16'b0100000000101100: out_v[126] = 10'b1100010111;
    16'b0000000000001000: out_v[126] = 10'b1011100101;
    16'b0000000000110000: out_v[126] = 10'b1001100101;
    16'b0100000000010100: out_v[126] = 10'b0110000011;
    16'b0100000000001000: out_v[126] = 10'b0100010101;
    16'b0000000000011010: out_v[126] = 10'b1100011011;
    16'b0100000000111010: out_v[126] = 10'b0110010101;
    16'b0100000000110100: out_v[126] = 10'b1001101111;
    16'b0000100000011010: out_v[126] = 10'b0000110111;
    16'b0100000000110110: out_v[126] = 10'b1000111011;
    16'b0100000000111000: out_v[126] = 10'b0111111111;
    16'b0100000000110000: out_v[126] = 10'b0100010011;
    16'b0100000000000000: out_v[126] = 10'b1011101001;
    16'b0000000000010100: out_v[126] = 10'b0111100100;
    16'b0100000000010010: out_v[126] = 10'b1101000011;
    16'b0100000000101000: out_v[126] = 10'b1111010111;
    16'b0100000000001100: out_v[126] = 10'b0111000011;
    16'b0000000000011000: out_v[126] = 10'b0101001110;
    16'b0100000000011100: out_v[126] = 10'b1111101000;
    16'b0000000000100000: out_v[126] = 10'b1000110111;
    16'b0100010000010110: out_v[126] = 10'b0110000001;
    16'b0000000000010010: out_v[126] = 10'b0010001000;
    16'b0000000000110010: out_v[126] = 10'b1001000010;
    16'b0100000000110010: out_v[126] = 10'b0011110111;
    16'b0100000000100100: out_v[126] = 10'b1010100101;
    16'b0100000000111100: out_v[126] = 10'b0011101011;
    16'b0000000000010110: out_v[126] = 10'b0011001101;
    16'b0100000000000100: out_v[126] = 10'b0011010010;
    16'b0100010000010100: out_v[126] = 10'b1100100111;
    16'b0100000000100000: out_v[126] = 10'b1110000111;
    16'b0000000000000000: out_v[126] = 10'b1100011111;
    16'b0100000000011000: out_v[126] = 10'b1110111011;
    16'b0000000000101000: out_v[126] = 10'b1011100101;
    16'b0000000000111000: out_v[126] = 10'b0001011001;
    16'b0000000000011100: out_v[126] = 10'b0101011101;
    16'b0000000000011110: out_v[126] = 10'b0010001011;
    16'b0000100000010010: out_v[126] = 10'b1011001000;
    16'b0000000000111010: out_v[126] = 10'b1010011001;
    16'b0100000000011110: out_v[126] = 10'b0011101110;
    16'b0100000000111110: out_v[126] = 10'b1000010101;
    16'b0000100000110010: out_v[126] = 10'b1000010011;
    16'b0000100000100010: out_v[126] = 10'b0111111001;
    16'b0000100000000010: out_v[126] = 10'b0011111011;
    16'b0000000000000010: out_v[126] = 10'b0010100110;
    16'b0000100000000000: out_v[126] = 10'b0100011010;
    16'b0000000000001010: out_v[126] = 10'b0101100010;
    16'b0000100000001000: out_v[126] = 10'b0111011000;
    16'b0000100000001010: out_v[126] = 10'b1101110000;
    16'b0000100000101010: out_v[126] = 10'b1000100101;
    16'b0000100000011000: out_v[126] = 10'b0011010101;
    16'b0100100000110000: out_v[126] = 10'b0111011100;
    16'b0000100000010000: out_v[126] = 10'b1101101010;
    16'b0000100000111010: out_v[126] = 10'b1111001101;
    16'b0100100000101000: out_v[126] = 10'b1111001111;
    16'b0000100000101000: out_v[126] = 10'b0111001110;
    16'b0100100000010000: out_v[126] = 10'b0110011010;
    16'b0000100000111000: out_v[126] = 10'b0111010000;
    16'b0000100000110000: out_v[126] = 10'b1011100100;
    16'b0000100000100000: out_v[126] = 10'b1000100110;
    16'b0000000000101010: out_v[126] = 10'b0001101010;
    16'b0000000000100010: out_v[126] = 10'b0111011000;
    16'b0000100000010110: out_v[126] = 10'b1101110100;
    16'b0000000000000100: out_v[126] = 10'b1000001011;
    16'b0100100000000100: out_v[126] = 10'b0000011001;
    16'b0000100000000110: out_v[126] = 10'b1000111010;
    16'b0000100000000100: out_v[126] = 10'b0001011011;
    16'b0000100000100100: out_v[126] = 10'b0101100101;
    16'b0000110000000100: out_v[126] = 10'b0101011011;
    16'b0000000000100100: out_v[126] = 10'b0000110101;
    16'b0000000000000110: out_v[126] = 10'b1010001011;
    16'b0100100000000000: out_v[126] = 10'b1110100001;
    16'b0100110000000100: out_v[126] = 10'b0110011011;
    16'b0000100000100110: out_v[126] = 10'b0111011000;
    16'b0000110000010110: out_v[126] = 10'b0100010101;
    16'b0000100000110110: out_v[126] = 10'b0111010110;
    16'b0100000000000010: out_v[126] = 10'b0111101010;
    16'b0100100000000010: out_v[126] = 10'b1100100111;
    16'b0000000000110100: out_v[126] = 10'b0011001011;
    16'b0000100000010100: out_v[126] = 10'b1101100111;
    16'b0000000000101100: out_v[126] = 10'b1001100010;
    16'b0000000000001100: out_v[126] = 10'b0001110010;
    16'b0001000000001000: out_v[126] = 10'b1010100010;
    16'b0001100000001000: out_v[126] = 10'b1101010011;
    16'b0100100000000110: out_v[126] = 10'b1011101110;
    16'b0100100000001000: out_v[126] = 10'b1110001111;
    16'b0000100000001100: out_v[126] = 10'b1001001011;
    16'b0000010000010110: out_v[126] = 10'b0110110111;
    16'b0000010000010000: out_v[126] = 10'b1000011100;
    16'b0000010000000110: out_v[126] = 10'b1100100101;
    16'b0000010000010010: out_v[126] = 10'b0100011111;
    16'b0100000000000110: out_v[126] = 10'b1111001011;
    16'b0100010000000110: out_v[126] = 10'b0111101000;
    16'b0000010000000010: out_v[126] = 10'b1100001011;
    16'b0100010000010010: out_v[126] = 10'b1101010010;
    16'b0100100000010010: out_v[126] = 10'b1110000010;
    16'b0100010000000010: out_v[126] = 10'b1100101001;
    16'b0100100000110010: out_v[126] = 10'b0101010000;
    16'b0100100000100000: out_v[126] = 10'b1010001100;
    16'b0100100000010100: out_v[126] = 10'b1000101101;
    16'b0100100000010110: out_v[126] = 10'b1100100011;
    default: out_v[126] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001001000000000: out_v[127] = 10'b1110100101;
    16'b0001000000000000: out_v[127] = 10'b0110001001;
    16'b0001000100000000: out_v[127] = 10'b0101100010;
    16'b0001010000000000: out_v[127] = 10'b1000101101;
    16'b0001100000000000: out_v[127] = 10'b0010011001;
    16'b0001110000000000: out_v[127] = 10'b0010010101;
    16'b0000010000000000: out_v[127] = 10'b1011101110;
    16'b0000011000000000: out_v[127] = 10'b1001001011;
    16'b0001010100000000: out_v[127] = 10'b1101011101;
    16'b0000000000000000: out_v[127] = 10'b0000011111;
    16'b0001011000000000: out_v[127] = 10'b0100000001;
    16'b0010011000000000: out_v[127] = 10'b0010101011;
    16'b0001100100000000: out_v[127] = 10'b1000100011;
    16'b0011011000000000: out_v[127] = 10'b0110111001;
    16'b0000100000000000: out_v[127] = 10'b0111010000;
    16'b0000001000000000: out_v[127] = 10'b0000101111;
    16'b0001111000000000: out_v[127] = 10'b1011011111;
    16'b0001101000000000: out_v[127] = 10'b1011011110;
    16'b0011101000000000: out_v[127] = 10'b0100110110;
    16'b0000101000000000: out_v[127] = 10'b0101000110;
    16'b0010001000000000: out_v[127] = 10'b1010001110;
    16'b0000110000000000: out_v[127] = 10'b1101010110;
    16'b0010101000000000: out_v[127] = 10'b0100011100;
    16'b0000111000000000: out_v[127] = 10'b1011010111;
    16'b0011001000000000: out_v[127] = 10'b1101100010;
    16'b0000100100000000: out_v[127] = 10'b0010110011;
    16'b0000000100000000: out_v[127] = 10'b1110101100;
    16'b0001001100000000: out_v[127] = 10'b0011100100;
    16'b0001100000001000: out_v[127] = 10'b1101100011;
    16'b0001100000100000: out_v[127] = 10'b1000001000;
    16'b0001000000100000: out_v[127] = 10'b1000101110;
    16'b0000100000100000: out_v[127] = 10'b1000110001;
    16'b0001100000000001: out_v[127] = 10'b1011101000;
    default: out_v[127] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100100010000101: out_v[128] = 10'b0100100001;
    16'b0100100110000101: out_v[128] = 10'b0000111011;
    16'b0100100110000000: out_v[128] = 10'b1000100011;
    16'b0100000010000101: out_v[128] = 10'b1001001011;
    16'b0100100010000000: out_v[128] = 10'b1010111001;
    16'b0100000010000100: out_v[128] = 10'b1000000101;
    16'b0100100010000001: out_v[128] = 10'b0110110100;
    16'b0100100100000101: out_v[128] = 10'b0101111101;
    16'b0100100010000100: out_v[128] = 10'b0001011100;
    16'b0100110110000000: out_v[128] = 10'b1011011011;
    16'b0100100000000101: out_v[128] = 10'b0100100111;
    16'b0100000110000100: out_v[128] = 10'b0011111001;
    16'b0000100010000001: out_v[128] = 10'b1001110101;
    16'b0100110110000101: out_v[128] = 10'b0001010001;
    16'b0101100110000100: out_v[128] = 10'b0111100101;
    16'b0100110110000100: out_v[128] = 10'b0001011100;
    16'b0100110010000101: out_v[128] = 10'b1010111101;
    16'b0100100110000100: out_v[128] = 10'b0110000101;
    16'b0100000010000001: out_v[128] = 10'b0010101010;
    16'b0100100110000001: out_v[128] = 10'b0011011001;
    16'b0100010110000100: out_v[128] = 10'b1111101000;
    16'b0100000000000101: out_v[128] = 10'b0101111011;
    16'b0100000110000000: out_v[128] = 10'b1001000011;
    16'b0000100010000000: out_v[128] = 10'b0110000111;
    16'b0100000000000001: out_v[128] = 10'b1001110001;
    16'b0100110010000100: out_v[128] = 10'b1011000110;
    16'b0000100110000000: out_v[128] = 10'b1110101100;
    16'b0000000010000101: out_v[128] = 10'b1001011001;
    16'b0000100010000101: out_v[128] = 10'b0101110001;
    16'b0100010110000000: out_v[128] = 10'b0011010011;
    16'b0100000010000000: out_v[128] = 10'b1000001010;
    16'b0000000000000000: out_v[128] = 10'b0101011101;
    16'b0000000010000000: out_v[128] = 10'b0101010011;
    16'b0000000000000001: out_v[128] = 10'b1010111101;
    16'b0000100000000001: out_v[128] = 10'b1001010111;
    16'b0100000000000000: out_v[128] = 10'b0110101110;
    16'b0100000000000100: out_v[128] = 10'b0000100110;
    16'b0000000010000001: out_v[128] = 10'b1111000010;
    16'b0000100000000000: out_v[128] = 10'b0011001111;
    16'b0000000000000100: out_v[128] = 10'b0010111110;
    16'b0100010010000000: out_v[128] = 10'b0111111010;
    16'b0100010011000100: out_v[128] = 10'b1010110101;
    16'b0100010010000100: out_v[128] = 10'b0010110011;
    16'b0100010000000100: out_v[128] = 10'b1111111011;
    16'b0000000010000100: out_v[128] = 10'b1110100001;
    16'b0000100000000100: out_v[128] = 10'b1000101110;
    16'b0100110000000100: out_v[128] = 10'b0111010011;
    16'b0000010000000100: out_v[128] = 10'b1110000111;
    16'b0100100000000100: out_v[128] = 10'b0011000100;
    16'b0100110010000000: out_v[128] = 10'b1010101011;
    16'b0100100000000000: out_v[128] = 10'b0111011000;
    16'b0100011001000100: out_v[128] = 10'b1100101101;
    16'b0100001010000000: out_v[128] = 10'b0011100110;
    16'b0100001010000100: out_v[128] = 10'b1001110110;
    16'b0100110001000100: out_v[128] = 10'b0110001001;
    16'b0100010001000100: out_v[128] = 10'b0101011010;
    16'b0000110001000100: out_v[128] = 10'b0001100111;
    16'b0000110000000100: out_v[128] = 10'b1000101111;
    16'b0100011011000100: out_v[128] = 10'b0110010111;
    16'b0100001000000100: out_v[128] = 10'b1100110110;
    16'b0100010011000000: out_v[128] = 10'b1011010100;
    16'b0100011011000000: out_v[128] = 10'b0100000011;
    16'b0000100000000101: out_v[128] = 10'b0110111000;
    16'b0100010000000000: out_v[128] = 10'b0111001111;
    16'b0000010001000100: out_v[128] = 10'b0011111111;
    16'b0100011010000100: out_v[128] = 10'b1100000111;
    16'b0000000000000101: out_v[128] = 10'b1000111001;
    16'b0100110011000100: out_v[128] = 10'b1011111111;
    16'b0000011010000001: out_v[128] = 10'b0010011010;
    16'b0100101010000001: out_v[128] = 10'b0110001000;
    16'b0100001010000001: out_v[128] = 10'b1011010010;
    16'b0100011010000001: out_v[128] = 10'b0110100011;
    16'b0100111010000001: out_v[128] = 10'b1011001110;
    16'b0000001010000001: out_v[128] = 10'b1100101100;
    16'b0100011010000000: out_v[128] = 10'b1011111100;
    16'b0000111010000001: out_v[128] = 10'b0001011110;
    16'b0000001010000000: out_v[128] = 10'b1111100011;
    16'b0100010010000001: out_v[128] = 10'b1000110111;
    16'b0100011010000101: out_v[128] = 10'b1101010010;
    16'b0100101010000000: out_v[128] = 10'b1110110001;
    16'b0000000100000000: out_v[128] = 10'b1000010101;
    16'b0001001100000000: out_v[128] = 10'b1101110011;
    16'b0000001000000000: out_v[128] = 10'b0001110111;
    16'b0000000110000000: out_v[128] = 10'b0011001011;
    16'b0000100100000000: out_v[128] = 10'b1110000111;
    16'b0000100010000100: out_v[128] = 10'b0111110000;
    16'b0001011100000000: out_v[128] = 10'b0001111110;
    16'b0000001100000000: out_v[128] = 10'b1001110010;
    16'b0000000100000100: out_v[128] = 10'b0011010110;
    16'b0001000100000000: out_v[128] = 10'b1010111010;
    16'b0000100110000001: out_v[128] = 10'b0111011011;
    16'b0100100000000001: out_v[128] = 10'b0100110010;
    16'b0100110010000001: out_v[128] = 10'b1000110110;
    16'b0100000100000100: out_v[128] = 10'b0110111000;
    16'b0000000100000001: out_v[128] = 10'b0011001110;
    16'b0001100100000001: out_v[128] = 10'b0011011101;
    16'b0000000110000001: out_v[128] = 10'b1100101011;
    16'b0001100000000001: out_v[128] = 10'b0101011110;
    16'b0100100010010000: out_v[128] = 10'b1101111101;
    16'b0001100000000000: out_v[128] = 10'b1010100101;
    16'b0001000100000001: out_v[128] = 10'b0110001011;
    16'b0000101010000000: out_v[128] = 10'b1111110011;
    16'b0001100010000000: out_v[128] = 10'b1101011101;
    16'b0001100100000000: out_v[128] = 10'b0011001010;
    16'b0001000110000001: out_v[128] = 10'b0111100011;
    16'b0001000010000001: out_v[128] = 10'b1011000101;
    16'b0001000000000001: out_v[128] = 10'b1011001111;
    16'b0001100110000001: out_v[128] = 10'b0011111100;
    16'b0001100110000000: out_v[128] = 10'b1001001100;
    16'b0100100010010001: out_v[128] = 10'b0011101111;
    16'b0001100010000001: out_v[128] = 10'b1000011100;
    16'b0000100100000001: out_v[128] = 10'b1101011101;
    16'b0000101000000000: out_v[128] = 10'b1101101001;
    16'b0101100010000000: out_v[128] = 10'b0001011110;
    16'b0100010010000101: out_v[128] = 10'b0101010010;
    16'b0000100100000100: out_v[128] = 10'b1101000111;
    16'b0001100100000100: out_v[128] = 10'b1000110111;
    16'b0000100100000101: out_v[128] = 10'b1000101101;
    16'b0001110100000000: out_v[128] = 10'b1100100110;
    default: out_v[128] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0101100001110000: out_v[129] = 10'b0011000011;
    16'b1100100001110000: out_v[129] = 10'b0001001111;
    16'b1101100001100000: out_v[129] = 10'b1111111100;
    16'b0101100001010000: out_v[129] = 10'b1011010011;
    16'b0101000001100000: out_v[129] = 10'b1001000100;
    16'b0101100001100000: out_v[129] = 10'b0101000100;
    16'b0001100000100000: out_v[129] = 10'b1000101110;
    16'b0001000000100000: out_v[129] = 10'b1100100101;
    16'b0101100001000000: out_v[129] = 10'b1001001011;
    16'b1100110001110000: out_v[129] = 10'b1100000011;
    16'b0101111001110000: out_v[129] = 10'b0111000100;
    16'b0100100001100000: out_v[129] = 10'b1101110111;
    16'b0100100001110000: out_v[129] = 10'b1110001111;
    16'b0100100001000000: out_v[129] = 10'b1000000100;
    16'b0101000000100000: out_v[129] = 10'b0011010011;
    16'b0101000001000000: out_v[129] = 10'b1001110111;
    16'b0001100001110000: out_v[129] = 10'b0011100111;
    16'b1101100001110000: out_v[129] = 10'b1111001001;
    16'b1100100001100000: out_v[129] = 10'b0001011001;
    16'b1101110001110000: out_v[129] = 10'b0000010011;
    16'b0001100001100000: out_v[129] = 10'b1101101000;
    16'b1100000001100000: out_v[129] = 10'b1000001010;
    16'b1101000001100000: out_v[129] = 10'b0001100100;
    16'b0101100001100010: out_v[129] = 10'b1101001011;
    16'b0100000001100000: out_v[129] = 10'b0101111110;
    16'b0101010001110000: out_v[129] = 10'b0011010101;
    16'b0101100000100000: out_v[129] = 10'b1000001110;
    16'b1100100001000000: out_v[129] = 10'b0011110011;
    16'b0001100001000000: out_v[129] = 10'b1111001011;
    16'b0101110001110000: out_v[129] = 10'b1000010001;
    16'b0101000001010000: out_v[129] = 10'b1101101001;
    16'b0100000001000000: out_v[129] = 10'b0001110111;
    16'b1101111001110000: out_v[129] = 10'b1010101111;
    16'b0101000001110000: out_v[129] = 10'b0100111011;
    16'b1001011001000000: out_v[129] = 10'b1001100011;
    16'b0001011001100000: out_v[129] = 10'b0000011011;
    16'b0100011000100000: out_v[129] = 10'b0111110111;
    16'b0000011000100000: out_v[129] = 10'b0101111001;
    16'b0000011001100000: out_v[129] = 10'b1101000011;
    16'b0100001000100000: out_v[129] = 10'b0111100111;
    16'b1001011001010000: out_v[129] = 10'b0001111100;
    16'b0100011000000000: out_v[129] = 10'b0100011011;
    16'b0001011001000000: out_v[129] = 10'b1001100011;
    16'b0001011001110000: out_v[129] = 10'b1101000111;
    16'b0100011000110000: out_v[129] = 10'b0110100011;
    16'b1001011000000000: out_v[129] = 10'b0101111111;
    16'b1001011001110000: out_v[129] = 10'b1001100011;
    16'b0000001000100000: out_v[129] = 10'b1000001111;
    16'b1001011001100000: out_v[129] = 10'b1111010001;
    16'b0001001001100000: out_v[129] = 10'b0110010101;
    16'b0001001001000000: out_v[129] = 10'b1000101110;
    16'b0101011001110000: out_v[129] = 10'b0011011110;
    16'b0100010000000000: out_v[129] = 10'b1111001011;
    16'b0101011001100000: out_v[129] = 10'b0000011100;
    16'b0100011001100000: out_v[129] = 10'b0001011001;
    16'b0000001001100000: out_v[129] = 10'b0111100010;
    16'b1001001001000000: out_v[129] = 10'b0010001011;
    16'b0000010000100000: out_v[129] = 10'b1110010110;
    16'b0101011001100010: out_v[129] = 10'b0111010111;
    16'b0101111001010000: out_v[129] = 10'b0111010110;
    16'b0101001001100000: out_v[129] = 10'b0010011100;
    16'b0101001001100010: out_v[129] = 10'b1111010010;
    16'b0001111000110000: out_v[129] = 10'b0101001011;
    16'b0101111000110000: out_v[129] = 10'b1101001000;
    16'b1001100001100000: out_v[129] = 10'b1011101011;
    16'b1101000001000000: out_v[129] = 10'b1011010101;
    16'b0001100000110000: out_v[129] = 10'b0111011110;
    16'b0001101000110000: out_v[129] = 10'b0001111111;
    16'b0001100000000000: out_v[129] = 10'b0111101101;
    16'b0101111001110010: out_v[129] = 10'b0000110111;
    16'b1101001001000000: out_v[129] = 10'b1111000101;
    16'b0001100000010000: out_v[129] = 10'b0110001101;
    16'b0001101000010000: out_v[129] = 10'b1011110010;
    16'b0001101000000000: out_v[129] = 10'b1001101001;
    16'b0101011001110010: out_v[129] = 10'b1111101011;
    16'b0001011000100000: out_v[129] = 10'b0101001010;
    16'b0000111000110000: out_v[129] = 10'b1010100110;
    16'b0101000001100010: out_v[129] = 10'b1111111010;
    16'b1101001001100000: out_v[129] = 10'b1001010111;
    16'b0101011001000000: out_v[129] = 10'b0100100011;
    16'b0001000001000000: out_v[129] = 10'b0010101100;
    16'b0001101000100000: out_v[129] = 10'b1001001010;
    16'b0001111001110000: out_v[129] = 10'b0111010110;
    16'b0101000001000010: out_v[129] = 10'b0011011111;
    16'b0001001000100000: out_v[129] = 10'b1100101111;
    16'b0001111000010000: out_v[129] = 10'b1000100101;
    16'b0001100001010000: out_v[129] = 10'b0010111011;
    16'b0101011001010000: out_v[129] = 10'b0110101010;
    16'b0101001001000000: out_v[129] = 10'b1001111010;
    16'b0001111001010000: out_v[129] = 10'b1110010010;
    16'b1001000001100000: out_v[129] = 10'b0010010000;
    16'b0101111000010000: out_v[129] = 10'b1011000111;
    16'b0101001001000010: out_v[129] = 10'b1111110000;
    16'b0000101000110000: out_v[129] = 10'b0110010101;
    16'b0101001000100000: out_v[129] = 10'b0000011110;
    16'b1100011001010000: out_v[129] = 10'b1011110010;
    16'b1100011001110000: out_v[129] = 10'b0010110111;
    16'b1101011001110000: out_v[129] = 10'b1011011010;
    16'b1100011001010010: out_v[129] = 10'b1111010111;
    16'b0000011001110010: out_v[129] = 10'b1111101010;
    16'b0100011001110010: out_v[129] = 10'b1011011000;
    16'b0100011001110000: out_v[129] = 10'b0011001010;
    16'b1100111001010000: out_v[129] = 10'b1100010110;
    16'b0000011000110000: out_v[129] = 10'b1011010101;
    16'b1101011001010000: out_v[129] = 10'b0011011011;
    16'b0000011001110000: out_v[129] = 10'b1001100101;
    16'b0100011000111000: out_v[129] = 10'b1001001110;
    16'b1100011001000000: out_v[129] = 10'b1100110100;
    16'b1101011001110010: out_v[129] = 10'b1000101011;
    16'b0100011001010000: out_v[129] = 10'b1011101011;
    16'b1100011001100000: out_v[129] = 10'b1110100001;
    16'b0100011001000000: out_v[129] = 10'b1101110101;
    16'b1100011001110010: out_v[129] = 10'b0110010110;
    16'b1100111001110000: out_v[129] = 10'b0101011010;
    16'b1101011001100000: out_v[129] = 10'b1101101001;
    16'b1101011001000000: out_v[129] = 10'b1111110011;
    16'b1100011001100010: out_v[129] = 10'b0101110111;
    16'b0100111001110000: out_v[129] = 10'b0100111010;
    16'b0000011001010000: out_v[129] = 10'b0000111001;
    16'b0000101000000000: out_v[129] = 10'b1001001101;
    16'b0000101000100000: out_v[129] = 10'b1110000010;
    16'b0100011000011000: out_v[129] = 10'b0010111111;
    16'b0000111001010000: out_v[129] = 10'b0100000110;
    16'b0000100000000010: out_v[129] = 10'b1100011100;
    16'b0000101001010000: out_v[129] = 10'b1000010010;
    16'b0100011000010000: out_v[129] = 10'b0101010101;
    16'b0100101000000000: out_v[129] = 10'b1100111011;
    16'b0100111000010000: out_v[129] = 10'b0000111110;
    16'b0100001000010000: out_v[129] = 10'b0101011001;
    16'b0000000000010000: out_v[129] = 10'b0001111011;
    16'b0000101001000000: out_v[129] = 10'b1001011001;
    16'b0000100000010000: out_v[129] = 10'b0100011001;
    16'b0100100000010000: out_v[129] = 10'b0101011010;
    16'b0000101000010000: out_v[129] = 10'b0111011001;
    16'b0100101000010000: out_v[129] = 10'b0111111100;
    16'b0100100000000000: out_v[129] = 10'b0100110010;
    16'b0000111000010000: out_v[129] = 10'b0011011000;
    16'b0100101000100000: out_v[129] = 10'b0111110011;
    16'b0000100000000000: out_v[129] = 10'b0110111000;
    16'b0000011000010000: out_v[129] = 10'b1010000011;
    16'b0000100000010010: out_v[129] = 10'b1010011010;
    16'b0000001000010000: out_v[129] = 10'b1101011011;
    16'b0100000000010000: out_v[129] = 10'b1101010010;
    16'b0100101000110000: out_v[129] = 10'b0110110000;
    16'b0100111000110000: out_v[129] = 10'b1010010011;
    16'b0000000000000000: out_v[129] = 10'b1010011110;
    16'b0100111000011000: out_v[129] = 10'b0101110011;
    16'b0000100000100000: out_v[129] = 10'b1001001110;
    16'b0001011001010000: out_v[129] = 10'b0101011000;
    16'b0100100000100000: out_v[129] = 10'b0011101110;
    16'b0100001000110000: out_v[129] = 10'b1111010101;
    16'b0000100000110000: out_v[129] = 10'b0011100111;
    16'b0100100000110000: out_v[129] = 10'b0111111010;
    16'b0100010001110000: out_v[129] = 10'b0010101000;
    16'b1100000001110000: out_v[129] = 10'b1111111100;
    16'b0101011101110001: out_v[129] = 10'b1100011100;
    16'b1100010001110000: out_v[129] = 10'b0011111110;
    16'b0001011000010000: out_v[129] = 10'b1010100111;
    16'b0001011000110000: out_v[129] = 10'b0100101000;
    16'b1100011101110001: out_v[129] = 10'b0111110101;
    16'b1100000101110001: out_v[129] = 10'b1111110110;
    16'b0101011000110000: out_v[129] = 10'b0010111011;
    16'b0100000001110000: out_v[129] = 10'b1010101110;
    16'b0001010000010000: out_v[129] = 10'b1110011000;
    16'b0101100000110000: out_v[129] = 10'b1000000111;
    16'b0101001000010000: out_v[129] = 10'b1111111010;
    16'b0101101000010000: out_v[129] = 10'b1011101111;
    16'b0101101000000000: out_v[129] = 10'b1000110111;
    16'b0101010000110000: out_v[129] = 10'b0010001101;
    16'b0101100000010000: out_v[129] = 10'b1010111101;
    16'b0101101000110000: out_v[129] = 10'b1010100111;
    16'b0100010000110000: out_v[129] = 10'b1101011001;
    16'b0101100000000000: out_v[129] = 10'b1011010001;
    16'b0101101001110000: out_v[129] = 10'b0000111011;
    16'b0101000000110000: out_v[129] = 10'b0000111111;
    16'b0101111000000000: out_v[129] = 10'b0101110100;
    16'b0101000000010000: out_v[129] = 10'b1110111011;
    16'b0101110000110000: out_v[129] = 10'b1101110100;
    16'b0101101000100000: out_v[129] = 10'b1111010010;
    16'b0100010000010000: out_v[129] = 10'b0011001001;
    16'b0101011000010000: out_v[129] = 10'b1110100000;
    16'b0101101001000000: out_v[129] = 10'b1011100001;
    16'b0001000001100000: out_v[129] = 10'b0010111001;
    16'b0100000000100000: out_v[129] = 10'b0011000111;
    16'b0100000000101000: out_v[129] = 10'b0111010010;
    16'b0100000010000000: out_v[129] = 10'b1101111001;
    16'b0000001001101000: out_v[129] = 10'b0111101101;
    16'b0000000001100000: out_v[129] = 10'b0111101000;
    16'b0100000010100000: out_v[129] = 10'b1110111010;
    16'b0000000000101000: out_v[129] = 10'b0001111101;
    16'b0100000001101000: out_v[129] = 10'b0111010010;
    16'b0100001000101000: out_v[129] = 10'b0101111011;
    16'b0100001010100000: out_v[129] = 10'b0111110001;
    16'b0100000000001000: out_v[129] = 10'b1000001111;
    16'b1001001001100000: out_v[129] = 10'b0011110011;
    16'b0001001001101000: out_v[129] = 10'b0011100101;
    16'b0100001001101000: out_v[129] = 10'b0011111001;
    16'b0100000000000000: out_v[129] = 10'b0011010000;
    16'b0000000010000000: out_v[129] = 10'b0010001111;
    16'b0000001000101000: out_v[129] = 10'b0011100000;
    16'b0100000000111000: out_v[129] = 10'b1011101111;
    16'b0000000001101000: out_v[129] = 10'b0101110011;
    16'b0000000000100000: out_v[129] = 10'b1011000001;
    16'b0000000010100000: out_v[129] = 10'b0111010011;
    16'b0100100000101000: out_v[129] = 10'b1100000100;
    16'b0100100010100000: out_v[129] = 10'b1010101110;
    16'b0101001001010000: out_v[129] = 10'b1101111011;
    16'b0101001001110000: out_v[129] = 10'b0110100011;
    16'b1000011001110000: out_v[129] = 10'b1111111101;
    16'b1000111001110000: out_v[129] = 10'b0111100110;
    16'b0101011001111000: out_v[129] = 10'b0101001111;
    16'b0100111001010000: out_v[129] = 10'b0100000110;
    16'b1001111001110000: out_v[129] = 10'b1000000111;
    16'b0001011001111000: out_v[129] = 10'b0110000011;
    16'b0100111001111000: out_v[129] = 10'b1111100001;
    16'b0000011000111000: out_v[129] = 10'b1011000100;
    16'b0100111000111000: out_v[129] = 10'b1011001000;
    16'b0100011001111000: out_v[129] = 10'b1001110111;
    16'b0100001000111000: out_v[129] = 10'b1110100011;
    16'b0100101000101000: out_v[129] = 10'b1001000111;
    16'b0000011001111000: out_v[129] = 10'b1001100111;
    16'b0000001000111000: out_v[129] = 10'b1001001111;
    16'b0100101010100000: out_v[129] = 10'b1101001010;
    16'b0100111010110000: out_v[129] = 10'b1000100010;
    16'b0100101000111000: out_v[129] = 10'b0101100110;
    16'b0000000000110000: out_v[129] = 10'b1001100110;
    16'b0000001000110000: out_v[129] = 10'b0100111100;
    16'b0100001010110000: out_v[129] = 10'b0100000111;
    16'b0000001001110000: out_v[129] = 10'b1100100111;
    16'b0100011010110000: out_v[129] = 10'b1000100001;
    16'b0100000000110000: out_v[129] = 10'b1000100111;
    default: out_v[129] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0111000000000000: out_v[130] = 10'b1101000101;
    16'b0110100011000100: out_v[130] = 10'b1100000110;
    16'b0100100011001110: out_v[130] = 10'b0111010111;
    16'b0100100001000110: out_v[130] = 10'b0010110001;
    16'b0111000000000100: out_v[130] = 10'b1001000011;
    16'b0110100000000100: out_v[130] = 10'b0001010110;
    16'b0100100000001110: out_v[130] = 10'b1111010011;
    16'b0010100010001100: out_v[130] = 10'b1110011011;
    16'b0100100011000110: out_v[130] = 10'b1011101011;
    16'b0100100010000110: out_v[130] = 10'b1011010100;
    16'b0110100011001100: out_v[130] = 10'b1011000111;
    16'b0000100000001110: out_v[130] = 10'b0101010011;
    16'b0010100010000100: out_v[130] = 10'b0100111110;
    16'b0110100001000110: out_v[130] = 10'b0100010110;
    16'b0110000001000100: out_v[130] = 10'b1001110011;
    16'b0100100000000110: out_v[130] = 10'b0111001011;
    16'b0111000001000100: out_v[130] = 10'b1111010001;
    16'b0110100000000110: out_v[130] = 10'b0111110110;
    16'b0110100001000100: out_v[130] = 10'b0011100110;
    16'b0111100000000110: out_v[130] = 10'b0011110011;
    16'b0000100010000110: out_v[130] = 10'b1101111100;
    16'b0110100001001100: out_v[130] = 10'b1111001010;
    16'b0100100001000010: out_v[130] = 10'b0111110010;
    16'b0101100000000110: out_v[130] = 10'b1001101001;
    16'b0110100011000110: out_v[130] = 10'b0011101011;
    16'b0111100001001100: out_v[130] = 10'b0011110101;
    16'b0100100000000010: out_v[130] = 10'b0110011001;
    16'b0100100000000100: out_v[130] = 10'b1101010011;
    16'b0000100000000110: out_v[130] = 10'b1001101010;
    16'b0100000000000110: out_v[130] = 10'b0010111010;
    16'b0000100001000010: out_v[130] = 10'b0001001111;
    16'b0111100000000100: out_v[130] = 10'b0001010110;
    16'b0100100001000100: out_v[130] = 10'b1101000111;
    16'b0110110011001100: out_v[130] = 10'b1101001111;
    16'b0101000000000100: out_v[130] = 10'b0111010101;
    16'b0111100000001110: out_v[130] = 10'b1001000011;
    16'b0110110011000100: out_v[130] = 10'b0111011111;
    16'b0111000001001100: out_v[130] = 10'b1011100101;
    16'b0100100001001110: out_v[130] = 10'b1101011111;
    16'b0000100000000010: out_v[130] = 10'b0010010011;
    16'b0110100011001110: out_v[130] = 10'b0001111110;
    16'b0111000000000110: out_v[130] = 10'b1111010011;
    16'b0110000000000100: out_v[130] = 10'b1000101001;
    16'b0111000000001100: out_v[130] = 10'b1001011001;
    16'b0001010001001000: out_v[130] = 10'b1010110111;
    16'b0000000000001100: out_v[130] = 10'b1100001011;
    16'b0100000000001100: out_v[130] = 10'b0000000011;
    16'b0100000000000100: out_v[130] = 10'b1110111001;
    16'b0000000000001000: out_v[130] = 10'b1000111011;
    16'b0000000001001000: out_v[130] = 10'b0001001111;
    16'b0000000000000000: out_v[130] = 10'b1101011011;
    16'b0001000001001000: out_v[130] = 10'b1110110010;
    16'b0000010001000000: out_v[130] = 10'b1111101001;
    16'b0001010000001000: out_v[130] = 10'b1011011011;
    16'b0001010000000000: out_v[130] = 10'b0110100011;
    16'b0000000000000100: out_v[130] = 10'b1101001110;
    16'b0001000001001100: out_v[130] = 10'b0000100011;
    16'b0000000001000000: out_v[130] = 10'b0111110001;
    16'b0001000011001000: out_v[130] = 10'b1111111101;
    16'b0000000001001100: out_v[130] = 10'b1001001110;
    16'b0101000000001100: out_v[130] = 10'b0110010010;
    16'b0000010001001000: out_v[130] = 10'b0111111101;
    16'b0001000010000000: out_v[130] = 10'b0011010110;
    16'b0001000000001000: out_v[130] = 10'b1000100111;
    16'b0001000000001100: out_v[130] = 10'b1011000101;
    16'b0001010001000000: out_v[130] = 10'b1001111011;
    16'b0000100000000100: out_v[130] = 10'b0101110001;
    16'b0100000001000100: out_v[130] = 10'b0101110101;
    16'b0001000000000000: out_v[130] = 10'b0010110100;
    16'b0000100000000000: out_v[130] = 10'b0001010111;
    16'b0000000001000100: out_v[130] = 10'b1111110100;
    16'b0001000000000100: out_v[130] = 10'b0011000100;
    16'b0001100000000100: out_v[130] = 10'b1101111011;
    16'b0001000000000110: out_v[130] = 10'b0011000100;
    16'b0001100000000000: out_v[130] = 10'b1001000000;
    16'b0011100000000000: out_v[130] = 10'b0100111110;
    16'b0010100000000000: out_v[130] = 10'b0010011101;
    16'b0001000001000100: out_v[130] = 10'b0100110110;
    16'b0001010010000000: out_v[130] = 10'b1010111101;
    16'b0000000000000010: out_v[130] = 10'b0111001010;
    16'b0001000000000010: out_v[130] = 10'b0001001111;
    16'b0001110010000000: out_v[130] = 10'b0101001011;
    16'b0101000001000100: out_v[130] = 10'b0101110101;
    16'b0000000000000110: out_v[130] = 10'b1011011000;
    16'b0001000000001010: out_v[130] = 10'b0011100100;
    16'b0101000001000110: out_v[130] = 10'b1001011101;
    16'b0101000000000110: out_v[130] = 10'b0110111111;
    16'b0001100010000000: out_v[130] = 10'b0110110011;
    16'b0001100000001000: out_v[130] = 10'b1000000110;
    16'b0100000001000110: out_v[130] = 10'b0000101110;
    16'b0000100010000000: out_v[130] = 10'b1101011011;
    16'b0010100000000100: out_v[130] = 10'b0010110111;
    16'b0110000001001100: out_v[130] = 10'b1001001110;
    16'b0110000011000100: out_v[130] = 10'b1010101111;
    16'b0010000000001000: out_v[130] = 10'b0111011001;
    16'b0100000001000000: out_v[130] = 10'b1101110010;
    16'b0000000000001010: out_v[130] = 10'b1000001100;
    16'b0110000000001000: out_v[130] = 10'b1101101100;
    16'b0110000001001000: out_v[130] = 10'b1111011001;
    16'b0100000001001100: out_v[130] = 10'b1001011111;
    16'b0100000001001000: out_v[130] = 10'b1011100101;
    16'b0110000000001100: out_v[130] = 10'b0111001011;
    16'b0100000000001110: out_v[130] = 10'b0011111111;
    16'b0110000001000000: out_v[130] = 10'b0111010111;
    16'b0010000001000000: out_v[130] = 10'b1011101011;
    16'b0100000001001110: out_v[130] = 10'b0111010010;
    16'b0010000000000000: out_v[130] = 10'b1011101101;
    16'b0110100000001100: out_v[130] = 10'b0110101011;
    16'b0100000000001000: out_v[130] = 10'b0001001010;
    16'b0100000000000000: out_v[130] = 10'b1101111001;
    16'b0100000011000100: out_v[130] = 10'b1001011111;
    16'b0000000001000010: out_v[130] = 10'b0010011011;
    16'b0110000001001110: out_v[130] = 10'b0101101101;
    16'b0100000001000010: out_v[130] = 10'b0011011110;
    16'b0110000000000000: out_v[130] = 10'b1110100100;
    16'b0010000001001000: out_v[130] = 10'b1010001101;
    16'b0110000000001110: out_v[130] = 10'b1100110010;
    16'b0011000000000010: out_v[130] = 10'b1111001110;
    16'b0110100010000100: out_v[130] = 10'b0110110111;
    16'b0011000000000000: out_v[130] = 10'b1100100011;
    16'b0001100000000010: out_v[130] = 10'b1001100011;
    16'b0001100010000010: out_v[130] = 10'b0000011001;
    16'b0010000000000010: out_v[130] = 10'b1101110110;
    16'b0010000000001010: out_v[130] = 10'b1101010001;
    16'b0110100010000110: out_v[130] = 10'b0011010010;
    16'b0010100000000010: out_v[130] = 10'b0101101110;
    16'b0011100000000010: out_v[130] = 10'b0010111000;
    16'b0010100011000000: out_v[130] = 10'b0111011111;
    16'b0000100010000010: out_v[130] = 10'b0000110000;
    16'b0110000000000110: out_v[130] = 10'b1100110000;
    16'b0010100010000000: out_v[130] = 10'b0011110110;
    16'b0111100010000100: out_v[130] = 10'b0110110110;
    16'b0011100010000000: out_v[130] = 10'b1010011000;
    16'b0011100000001000: out_v[130] = 10'b1010001111;
    16'b0011100010000100: out_v[130] = 10'b0110001010;
    16'b0011000000001000: out_v[130] = 10'b0010110011;
    16'b0001110000000010: out_v[130] = 10'b1110011001;
    16'b0010000000000100: out_v[130] = 10'b0101101001;
    16'b0101100010000110: out_v[130] = 10'b1000110101;
    16'b0111100010000110: out_v[130] = 10'b1111011110;
    16'b0010100000001000: out_v[130] = 10'b0011011001;
    16'b0110000011000010: out_v[130] = 10'b0011010111;
    16'b0110000010000100: out_v[130] = 10'b1000111010;
    16'b0010000000001100: out_v[130] = 10'b0110001010;
    16'b0010000010000100: out_v[130] = 10'b1101110100;
    16'b0110000001000110: out_v[130] = 10'b1101110101;
    16'b0110000011000110: out_v[130] = 10'b1101010011;
    16'b0000000010000100: out_v[130] = 10'b1111001001;
    16'b0010000010000000: out_v[130] = 10'b1000100010;
    16'b0110000011001100: out_v[130] = 10'b1001101110;
    16'b0110010001000100: out_v[130] = 10'b1010111011;
    16'b0110000010000110: out_v[130] = 10'b1011001001;
    16'b0010000010001100: out_v[130] = 10'b1100110110;
    16'b0110000011000000: out_v[130] = 10'b1011011111;
    16'b0110000010001100: out_v[130] = 10'b1010110111;
    16'b0000000010001100: out_v[130] = 10'b0010110100;
    16'b0010000010001000: out_v[130] = 10'b1001100110;
    16'b0110010000000110: out_v[130] = 10'b1110111110;
    16'b0100000010000100: out_v[130] = 10'b1010100001;
    16'b0110010000000100: out_v[130] = 10'b0110111111;
    16'b0110000000000010: out_v[130] = 10'b1001110001;
    16'b0011100000000100: out_v[130] = 10'b1110011110;
    16'b0011000000001100: out_v[130] = 10'b1100000101;
    16'b0011000000010100: out_v[130] = 10'b1000100011;
    16'b0011110000000100: out_v[130] = 10'b1111110010;
    16'b0000100000010110: out_v[130] = 10'b0110111100;
    16'b0011000000000100: out_v[130] = 10'b0001011001;
    16'b0111010000000100: out_v[130] = 10'b1001011011;
    16'b0011100000000110: out_v[130] = 10'b1101111011;
    16'b0001100000000110: out_v[130] = 10'b0101010111;
    16'b0001100000010110: out_v[130] = 10'b1101011011;
    16'b0011010000000100: out_v[130] = 10'b1111000010;
    16'b0011100000010100: out_v[130] = 10'b0110111001;
    16'b0011010000001100: out_v[130] = 10'b1100001110;
    16'b0010000000010100: out_v[130] = 10'b1011001010;
    16'b0001000000010100: out_v[130] = 10'b1001000000;
    16'b0101010000001100: out_v[130] = 10'b1001011011;
    16'b0001010000001100: out_v[130] = 10'b1111001000;
    16'b0010100000010100: out_v[130] = 10'b1011011110;
    16'b0011000000000110: out_v[130] = 10'b1011101011;
    16'b0111010000001100: out_v[130] = 10'b0100101111;
    16'b0011000000010000: out_v[130] = 10'b0111001011;
    16'b0011100000010110: out_v[130] = 10'b1110110101;
    16'b0010110000000100: out_v[130] = 10'b1011001111;
    16'b0100000011001110: out_v[130] = 10'b0011001110;
    16'b0000000000001011: out_v[130] = 10'b0010011011;
    16'b0000100000001010: out_v[130] = 10'b0110001100;
    16'b0100000000101110: out_v[130] = 10'b0000111100;
    16'b0000000011000000: out_v[130] = 10'b0101111110;
    16'b0000000011000110: out_v[130] = 10'b0011101011;
    16'b0000000000001110: out_v[130] = 10'b0101010111;
    16'b0000000001000110: out_v[130] = 10'b0010110000;
    16'b0101000000001110: out_v[130] = 10'b0011101011;
    16'b0100000010001110: out_v[130] = 10'b1011000011;
    16'b0000000001001110: out_v[130] = 10'b0111111110;
    16'b0100000010000110: out_v[130] = 10'b1111100000;
    16'b0000000011001110: out_v[130] = 10'b1001010110;
    16'b0101000001000000: out_v[130] = 10'b1001010110;
    16'b0101000011000100: out_v[130] = 10'b1001111110;
    16'b0001000001000000: out_v[130] = 10'b0011001110;
    16'b0111000011000100: out_v[130] = 10'b0011111000;
    16'b0111000010000110: out_v[130] = 10'b1110000111;
    16'b0101000011000000: out_v[130] = 10'b1111011111;
    16'b0101000001001100: out_v[130] = 10'b0000010111;
    16'b0111000011000110: out_v[130] = 10'b0101010011;
    16'b0001000011000100: out_v[130] = 10'b0111010111;
    16'b0101010011000100: out_v[130] = 10'b0010010100;
    16'b0111000011000010: out_v[130] = 10'b1100110011;
    16'b0101000000000000: out_v[130] = 10'b0101001010;
    16'b0111000000001110: out_v[130] = 10'b1110110011;
    16'b0101000010000100: out_v[130] = 10'b1100100110;
    16'b0101000011001100: out_v[130] = 10'b1100110101;
    16'b0111000001000110: out_v[130] = 10'b0111100111;
    16'b0001000011000000: out_v[130] = 10'b1011101011;
    16'b0111000000000010: out_v[130] = 10'b0111000010;
    16'b0010000001000100: out_v[130] = 10'b1101100001;
    16'b0101100000000100: out_v[130] = 10'b1111001110;
    16'b0001100000001011: out_v[130] = 10'b1101011011;
    16'b0001100000001010: out_v[130] = 10'b1000111010;
    16'b0001100000000011: out_v[130] = 10'b1101001011;
    default: out_v[130] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000010011000: out_v[131] = 10'b0010100001;
    16'b0000000010001000: out_v[131] = 10'b1110100010;
    16'b0010000010001001: out_v[131] = 10'b0101001111;
    16'b0010000010001010: out_v[131] = 10'b1001010110;
    16'b0000000010011010: out_v[131] = 10'b1110010111;
    16'b1000000010101000: out_v[131] = 10'b1001000010;
    16'b0010001000000000: out_v[131] = 10'b1000110011;
    16'b0010000000001010: out_v[131] = 10'b0001100111;
    16'b0010001000001000: out_v[131] = 10'b0010011001;
    16'b0010000010001000: out_v[131] = 10'b1111100100;
    16'b1000000010111010: out_v[131] = 10'b0111001011;
    16'b0000000010000000: out_v[131] = 10'b0110001011;
    16'b1000000010001000: out_v[131] = 10'b1011100110;
    16'b0010000010000010: out_v[131] = 10'b0100101010;
    16'b1000000010011000: out_v[131] = 10'b1000111000;
    16'b1000000010001010: out_v[131] = 10'b0011011111;
    16'b0000000010001010: out_v[131] = 10'b0110001001;
    16'b0000000010001001: out_v[131] = 10'b0011101000;
    16'b0000000010010000: out_v[131] = 10'b1001001011;
    16'b0010000000001000: out_v[131] = 10'b1110000011;
    16'b0010001010001000: out_v[131] = 10'b1101110111;
    16'b1000000010101010: out_v[131] = 10'b0100000101;
    16'b0000000010000010: out_v[131] = 10'b1001110010;
    16'b0000000000001010: out_v[131] = 10'b1110011100;
    16'b0010000000000000: out_v[131] = 10'b0010110000;
    16'b1010000010101000: out_v[131] = 10'b1001101011;
    16'b0010000010101000: out_v[131] = 10'b0001001011;
    16'b1000000010111000: out_v[131] = 10'b1000001100;
    16'b0010001000001001: out_v[131] = 10'b0110100101;
    16'b1000000010011010: out_v[131] = 10'b0000111111;
    16'b0010000010011000: out_v[131] = 10'b1010011011;
    16'b0010000000000010: out_v[131] = 10'b1110001111;
    16'b0000000000001000: out_v[131] = 10'b1010100111;
    16'b1000000000111000: out_v[131] = 10'b1000110110;
    16'b0010001000001010: out_v[131] = 10'b1011110111;
    16'b0000000000011000: out_v[131] = 10'b0110101100;
    16'b0000000000111000: out_v[131] = 10'b0111101100;
    16'b0000000000100000: out_v[131] = 10'b0100111010;
    16'b0000000000000000: out_v[131] = 10'b1000110110;
    16'b0000000000100010: out_v[131] = 10'b1110000010;
    16'b0000000000010000: out_v[131] = 10'b0010110110;
    16'b0000000000000010: out_v[131] = 10'b1011010110;
    16'b1000000000100000: out_v[131] = 10'b0110010101;
    16'b1000000000111010: out_v[131] = 10'b0000110111;
    16'b0000000000110010: out_v[131] = 10'b1111001001;
    16'b1000000000100010: out_v[131] = 10'b1100110110;
    16'b0000000000010010: out_v[131] = 10'b1010011110;
    16'b0000000000101000: out_v[131] = 10'b0111101100;
    16'b0000000000111010: out_v[131] = 10'b1010101010;
    16'b0000000000011010: out_v[131] = 10'b1010110100;
    16'b0000000000110000: out_v[131] = 10'b1100101010;
    16'b0000000000101010: out_v[131] = 10'b1110010001;
    16'b1000000000111001: out_v[131] = 10'b0011011000;
    16'b0000000000010001: out_v[131] = 10'b1001110110;
    16'b1000000000101010: out_v[131] = 10'b0111011100;
    16'b1000000000110001: out_v[131] = 10'b0010111011;
    16'b1100000010110010: out_v[131] = 10'b0010100110;
    16'b1100000000111010: out_v[131] = 10'b0010101111;
    16'b1000000000110010: out_v[131] = 10'b0111011001;
    16'b1000000010110010: out_v[131] = 10'b1101001000;
    16'b1000000000110000: out_v[131] = 10'b1000011101;
    16'b0000000000011011: out_v[131] = 10'b1110011110;
    16'b1000000000101011: out_v[131] = 10'b1110111111;
    16'b1100000000110010: out_v[131] = 10'b1110001111;
    16'b1000000000101000: out_v[131] = 10'b0010001010;
    16'b1000000000111011: out_v[131] = 10'b0101110101;
    16'b1000000010110001: out_v[131] = 10'b0110000110;
    16'b0000000000011001: out_v[131] = 10'b1000110110;
    16'b1000000010110000: out_v[131] = 10'b0010011100;
    16'b1000000000011010: out_v[131] = 10'b0101110010;
    16'b1100000010111010: out_v[131] = 10'b1100010100;
    16'b0000000000110001: out_v[131] = 10'b0100001000;
    16'b1000000010100010: out_v[131] = 10'b0111100100;
    16'b1000000010111001: out_v[131] = 10'b0011111010;
    16'b1000000000101001: out_v[131] = 10'b1010000010;
    16'b1000000000100001: out_v[131] = 10'b0110110100;
    16'b0000001000110000: out_v[131] = 10'b1100101100;
    16'b1000000010001001: out_v[131] = 10'b0001100010;
    16'b1000000000000000: out_v[131] = 10'b1110001000;
    16'b1000000010011001: out_v[131] = 10'b0111011000;
    16'b1000000000001000: out_v[131] = 10'b0100111000;
    16'b1000000000001001: out_v[131] = 10'b0110011111;
    16'b1000000000010000: out_v[131] = 10'b1100101001;
    16'b1000000010000001: out_v[131] = 10'b1100011000;
    16'b1000000000000001: out_v[131] = 10'b1011001001;
    16'b1000000000000010: out_v[131] = 10'b0010101000;
    16'b1000000010000010: out_v[131] = 10'b0000100100;
    16'b0000000010000001: out_v[131] = 10'b0010011001;
    16'b1000000000011000: out_v[131] = 10'b1101001010;
    16'b1000000010000000: out_v[131] = 10'b0110011011;
    16'b1000000000001010: out_v[131] = 10'b0000001011;
    16'b1000000000010001: out_v[131] = 10'b0100011101;
    16'b1000000010010001: out_v[131] = 10'b1101010100;
    16'b1000000000011001: out_v[131] = 10'b1101000010;
    16'b1000000010100000: out_v[131] = 10'b0010010110;
    16'b1000000010010000: out_v[131] = 10'b1110010011;
    16'b1000001010111000: out_v[131] = 10'b1010000111;
    16'b1000001010110000: out_v[131] = 10'b0011101110;
    16'b1010000010110000: out_v[131] = 10'b0100010010;
    16'b1100000000010010: out_v[131] = 10'b1010111100;
    16'b1000000010010010: out_v[131] = 10'b1001011100;
    16'b1100000010010010: out_v[131] = 10'b1000001101;
    16'b1100000000111000: out_v[131] = 10'b0101010010;
    16'b1100000010100010: out_v[131] = 10'b0111001111;
    16'b1100000010111000: out_v[131] = 10'b0111110010;
    16'b1000000000010010: out_v[131] = 10'b0111010101;
    16'b1100000000011000: out_v[131] = 10'b1001011101;
    16'b0100000010010010: out_v[131] = 10'b0011001100;
    16'b0000000010010010: out_v[131] = 10'b1011100010;
    16'b0000000010110000: out_v[131] = 10'b0111000100;
    16'b1100000000110000: out_v[131] = 10'b0011010100;
    16'b0000000010100000: out_v[131] = 10'b1101001010;
    16'b0100000000110010: out_v[131] = 10'b1111011001;
    16'b1100000000010000: out_v[131] = 10'b0010111011;
    16'b1100000010010000: out_v[131] = 10'b1011111011;
    16'b1000000010101001: out_v[131] = 10'b0000000110;
    16'b1000000010100001: out_v[131] = 10'b1010001111;
    16'b1010000010111000: out_v[131] = 10'b1110001010;
    default: out_v[131] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1010000100001000: out_v[132] = 10'b1111000001;
    16'b0010000100001001: out_v[132] = 10'b1010100111;
    16'b1010000100011010: out_v[132] = 10'b0111001001;
    16'b1100000100001000: out_v[132] = 10'b0001010001;
    16'b1010000100000011: out_v[132] = 10'b0000111100;
    16'b1100000100011010: out_v[132] = 10'b1101000100;
    16'b1010000100001001: out_v[132] = 10'b0011001011;
    16'b1010000100001010: out_v[132] = 10'b1111100111;
    16'b1100000100001010: out_v[132] = 10'b1100101110;
    16'b0010000000001010: out_v[132] = 10'b1110100011;
    16'b0010000000000010: out_v[132] = 10'b0100111101;
    16'b0010000100001010: out_v[132] = 10'b1101101010;
    16'b1010000000001010: out_v[132] = 10'b1001110110;
    16'b1110000100001011: out_v[132] = 10'b1101001011;
    16'b1010000000000011: out_v[132] = 10'b0111111010;
    16'b1010000100000010: out_v[132] = 10'b0000110010;
    16'b1010001100001010: out_v[132] = 10'b1011100110;
    16'b1010000001000011: out_v[132] = 10'b0111000010;
    16'b1010000000000000: out_v[132] = 10'b1101101110;
    16'b1100000100001001: out_v[132] = 10'b0110100110;
    16'b1110000100001010: out_v[132] = 10'b0000011110;
    16'b1010000101000011: out_v[132] = 10'b0011001111;
    16'b1010000100001011: out_v[132] = 10'b1110100000;
    16'b1010000000011010: out_v[132] = 10'b1011001011;
    16'b1110000100001000: out_v[132] = 10'b1101110011;
    16'b1110000100011011: out_v[132] = 10'b1100010111;
    16'b0110000100001001: out_v[132] = 10'b1110011001;
    16'b1110000100001001: out_v[132] = 10'b0001111110;
    16'b0010000101000011: out_v[132] = 10'b1101110101;
    16'b1000000100001010: out_v[132] = 10'b0110001010;
    16'b0010000100001011: out_v[132] = 10'b0011111011;
    16'b0110000100011010: out_v[132] = 10'b1110110110;
    16'b1010000000000010: out_v[132] = 10'b0010011001;
    16'b1110000100011010: out_v[132] = 10'b0001100111;
    16'b1100000100011000: out_v[132] = 10'b1001011001;
    16'b0000000000000010: out_v[132] = 10'b0110011000;
    16'b0110000100011001: out_v[132] = 10'b0111001010;
    16'b0010000100000011: out_v[132] = 10'b0101110110;
    16'b0010000000011010: out_v[132] = 10'b1011000101;
    16'b0100000100011010: out_v[132] = 10'b0000110101;
    16'b1000000000000010: out_v[132] = 10'b1011001011;
    16'b0010000100011010: out_v[132] = 10'b1000011011;
    16'b1000000000010000: out_v[132] = 10'b1110110100;
    16'b0000000000000000: out_v[132] = 10'b0101010010;
    16'b0000000100000000: out_v[132] = 10'b1010001100;
    16'b0000000100000010: out_v[132] = 10'b1001010110;
    16'b0000000000010000: out_v[132] = 10'b1101100110;
    16'b1000000000000000: out_v[132] = 10'b1101101011;
    16'b0100000100000010: out_v[132] = 10'b0000011010;
    16'b1100000000010000: out_v[132] = 10'b1101000111;
    16'b1000000100010000: out_v[132] = 10'b0111001110;
    16'b0000000100010000: out_v[132] = 10'b0110011111;
    16'b0000001100000010: out_v[132] = 10'b0111001110;
    16'b1000000100000000: out_v[132] = 10'b1001110111;
    16'b0000000100010010: out_v[132] = 10'b0110110111;
    16'b0000000000010010: out_v[132] = 10'b0111110101;
    16'b0100000000010010: out_v[132] = 10'b0010000011;
    16'b1000000000010010: out_v[132] = 10'b1011110100;
    16'b1100000000011000: out_v[132] = 10'b0000111100;
    16'b1100000000000010: out_v[132] = 10'b0001011111;
    16'b1000000000010001: out_v[132] = 10'b1111110100;
    16'b0100000000010000: out_v[132] = 10'b0010110110;
    16'b1100000000001010: out_v[132] = 10'b0100101111;
    16'b0100000000011010: out_v[132] = 10'b0000101111;
    16'b0100000000011000: out_v[132] = 10'b0011001000;
    16'b1100000000011010: out_v[132] = 10'b1101001010;
    16'b1100000000010011: out_v[132] = 10'b0011110011;
    16'b0100000000001000: out_v[132] = 10'b0000110101;
    16'b1100000000011001: out_v[132] = 10'b1111111001;
    16'b1110000000011011: out_v[132] = 10'b1001111010;
    16'b1110000000011010: out_v[132] = 10'b1000111010;
    16'b1100000000011111: out_v[132] = 10'b1110011011;
    16'b1100000000010010: out_v[132] = 10'b0110001010;
    16'b0100000100010010: out_v[132] = 10'b0111100011;
    16'b1100000100011011: out_v[132] = 10'b1100101011;
    16'b1100000000001011: out_v[132] = 10'b1111011100;
    16'b1100000000011011: out_v[132] = 10'b0101100011;
    16'b1100000100010010: out_v[132] = 10'b0100000011;
    16'b1000000100010010: out_v[132] = 10'b1010111001;
    16'b1000000000011010: out_v[132] = 10'b0111001011;
    16'b1000000000010011: out_v[132] = 10'b0011110100;
    16'b1100000000010001: out_v[132] = 10'b0011001100;
    16'b0100000000001010: out_v[132] = 10'b1000000111;
    16'b1000000000011011: out_v[132] = 10'b1011100111;
    16'b1100000100010011: out_v[132] = 10'b0111010101;
    16'b1100000000001000: out_v[132] = 10'b0101111011;
    16'b1100000000001001: out_v[132] = 10'b0111110010;
    16'b1110000000001011: out_v[132] = 10'b1010010100;
    16'b0110000000011010: out_v[132] = 10'b1111000010;
    16'b0110000000010010: out_v[132] = 10'b1110100011;
    16'b0100000000000010: out_v[132] = 10'b1111100000;
    16'b1100000000011101: out_v[132] = 10'b0100011101;
    16'b0000000000011010: out_v[132] = 10'b0011010111;
    16'b1110000000011001: out_v[132] = 10'b1010111110;
    16'b1100000000000000: out_v[132] = 10'b1100011010;
    16'b1000000000011000: out_v[132] = 10'b0000001101;
    16'b0100000000000000: out_v[132] = 10'b1011101000;
    16'b0000000000001010: out_v[132] = 10'b1000001111;
    16'b0100001000000010: out_v[132] = 10'b1011001001;
    16'b1100001000000010: out_v[132] = 10'b1111001011;
    16'b1100000000000011: out_v[132] = 10'b0011011011;
    16'b0100001000001010: out_v[132] = 10'b1001000001;
    16'b0100001100000010: out_v[132] = 10'b0101111110;
    16'b1100000100000000: out_v[132] = 10'b1010001000;
    16'b1100000100000011: out_v[132] = 10'b1001001100;
    16'b0010001100000010: out_v[132] = 10'b0101110110;
    16'b1100000100000010: out_v[132] = 10'b1000100100;
    16'b1100001000001010: out_v[132] = 10'b1110000111;
    16'b1100000100001011: out_v[132] = 10'b0100001101;
    16'b1100000100000001: out_v[132] = 10'b1011001010;
    16'b0010000100000010: out_v[132] = 10'b1100001001;
    16'b1010000100000001: out_v[132] = 10'b1010001111;
    16'b1100000000000001: out_v[132] = 10'b1111000111;
    16'b0100000100001010: out_v[132] = 10'b0011001110;
    16'b0010000100000000: out_v[132] = 10'b0010100001;
    16'b1010000100000000: out_v[132] = 10'b1010111011;
    16'b1110000000001010: out_v[132] = 10'b0011111101;
    16'b1110000100000011: out_v[132] = 10'b0100011111;
    16'b1010000000001011: out_v[132] = 10'b0111011010;
    16'b1000000000001010: out_v[132] = 10'b1111000111;
    16'b1000000000000011: out_v[132] = 10'b1001011010;
    16'b0100000100000000: out_v[132] = 10'b1101001000;
    16'b1100001000011000: out_v[132] = 10'b0011111111;
    16'b0100000100001000: out_v[132] = 10'b1101101110;
    16'b1100001000001000: out_v[132] = 10'b0111000111;
    16'b0110000100001010: out_v[132] = 10'b0000111011;
    16'b0100001100001010: out_v[132] = 10'b0110010100;
    16'b0110000000001010: out_v[132] = 10'b0110010000;
    16'b1110000000011000: out_v[132] = 10'b0000011010;
    16'b0110000000001000: out_v[132] = 10'b1100110111;
    16'b0110001000001000: out_v[132] = 10'b1101111111;
    16'b0100001000001000: out_v[132] = 10'b0101111111;
    16'b1110000000001000: out_v[132] = 10'b1000110100;
    16'b0000000100011000: out_v[132] = 10'b1001111100;
    16'b0110000100011000: out_v[132] = 10'b1000011101;
    16'b0100000100011000: out_v[132] = 10'b1001001000;
    16'b0100001100011010: out_v[132] = 10'b1101100010;
    16'b0110000000011000: out_v[132] = 10'b0001110010;
    16'b0110000100001000: out_v[132] = 10'b1110001110;
    16'b0100001000011010: out_v[132] = 10'b1000101010;
    16'b0100001000000000: out_v[132] = 10'b0011010111;
    16'b0000000100001010: out_v[132] = 10'b1011010111;
    16'b1110000100011000: out_v[132] = 10'b1101110010;
    16'b0000000100001000: out_v[132] = 10'b1110101010;
    16'b0000000000001000: out_v[132] = 10'b0111111011;
    16'b0110000001001000: out_v[132] = 10'b0110011011;
    16'b0100001000011000: out_v[132] = 10'b0000111001;
    16'b0100000100000011: out_v[132] = 10'b1101110010;
    16'b1000000100000010: out_v[132] = 10'b1000110001;
    16'b0000000100001001: out_v[132] = 10'b1101110110;
    16'b0000000100011010: out_v[132] = 10'b1000111001;
    16'b0100000100010000: out_v[132] = 10'b1111101000;
    16'b0100000100001011: out_v[132] = 10'b1001110010;
    16'b0000000000011000: out_v[132] = 10'b0111101000;
    16'b1010001000001010: out_v[132] = 10'b1001100101;
    16'b0100000100000001: out_v[132] = 10'b1001110110;
    16'b0000000100000001: out_v[132] = 10'b0001001011;
    16'b0100000100001001: out_v[132] = 10'b1110100011;
    16'b1100001100001010: out_v[132] = 10'b1000110100;
    16'b1110000100011110: out_v[132] = 10'b1110111111;
    16'b1100000100010000: out_v[132] = 10'b0111001110;
    16'b1100000100001100: out_v[132] = 10'b0100000111;
    16'b1100000100011110: out_v[132] = 10'b0011011110;
    16'b0010000100010010: out_v[132] = 10'b1100101011;
    16'b1000000100011000: out_v[132] = 10'b0111011110;
    16'b0110000100010010: out_v[132] = 10'b1011011100;
    16'b1100000100011100: out_v[132] = 10'b0111101110;
    16'b1000000100011100: out_v[132] = 10'b1111111001;
    16'b1100000100010100: out_v[132] = 10'b1010111111;
    16'b1000000100011010: out_v[132] = 10'b0011010100;
    16'b0010000000010010: out_v[132] = 10'b1111110010;
    16'b0010000000011000: out_v[132] = 10'b0011000011;
    16'b1010000100011000: out_v[132] = 10'b0101111000;
    16'b1010000100011110: out_v[132] = 10'b0111011111;
    16'b1110000100011100: out_v[132] = 10'b0111001110;
    16'b1010000100011100: out_v[132] = 10'b0101111011;
    16'b0100001100000000: out_v[132] = 10'b1000011011;
    16'b0100001100001000: out_v[132] = 10'b1100001000;
    16'b0110000100000010: out_v[132] = 10'b0101001010;
    16'b0110000100000000: out_v[132] = 10'b0110000000;
    16'b0110000000000010: out_v[132] = 10'b1010101001;
    16'b1100001000010010: out_v[132] = 10'b1101001011;
    16'b1000001100010010: out_v[132] = 10'b0011010111;
    16'b0100001000010010: out_v[132] = 10'b1011010010;
    16'b1000001000010010: out_v[132] = 10'b1011010111;
    16'b1100001000011010: out_v[132] = 10'b0110011010;
    16'b0100001100010010: out_v[132] = 10'b0110110000;
    16'b1100001100010010: out_v[132] = 10'b1011001110;
    16'b1100001100011010: out_v[132] = 10'b1110101001;
    16'b1000000100010011: out_v[132] = 10'b1001111111;
    16'b0100000010001010: out_v[132] = 10'b1111100111;
    16'b0100001010001010: out_v[132] = 10'b1000001111;
    default: out_v[132] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1010010000001100: out_v[133] = 10'b0010101011;
    16'b0000110000111100: out_v[133] = 10'b1010111111;
    16'b1000010001101100: out_v[133] = 10'b0110100001;
    16'b1010010000101100: out_v[133] = 10'b0010110011;
    16'b0000010000100100: out_v[133] = 10'b0011001011;
    16'b0000110000011100: out_v[133] = 10'b0000110111;
    16'b0000010000101100: out_v[133] = 10'b0110100110;
    16'b0010010000001100: out_v[133] = 10'b1010110101;
    16'b1000010000101100: out_v[133] = 10'b0101110010;
    16'b0010110000111100: out_v[133] = 10'b0011000111;
    16'b0010110000001000: out_v[133] = 10'b0010100111;
    16'b0000110000101100: out_v[133] = 10'b0101010111;
    16'b0000100000110000: out_v[133] = 10'b1111100011;
    16'b0000110000101000: out_v[133] = 10'b1010111110;
    16'b0000110001011100: out_v[133] = 10'b0100101011;
    16'b0010100100110000: out_v[133] = 10'b1101001110;
    16'b0000110000111000: out_v[133] = 10'b1110101100;
    16'b0000010000111100: out_v[133] = 10'b1111010010;
    16'b0010100100110001: out_v[133] = 10'b1011110001;
    16'b1000010000100000: out_v[133] = 10'b1001011101;
    16'b1000110000101100: out_v[133] = 10'b1101001111;
    16'b0000110001111100: out_v[133] = 10'b1101011111;
    16'b1000010001000000: out_v[133] = 10'b1000100011;
    16'b0000110001101100: out_v[133] = 10'b0001110110;
    16'b0010110000011000: out_v[133] = 10'b0010001100;
    16'b0000100000111000: out_v[133] = 10'b0010010011;
    16'b0010110000011100: out_v[133] = 10'b0110110110;
    16'b0010100000010000: out_v[133] = 10'b1100010101;
    16'b1000000000100000: out_v[133] = 10'b0111110011;
    16'b0010110000001100: out_v[133] = 10'b1001000111;
    16'b1000110001101100: out_v[133] = 10'b1101011000;
    16'b0000010000101000: out_v[133] = 10'b1101000011;
    16'b0010100100010000: out_v[133] = 10'b0100110011;
    16'b1000010000001100: out_v[133] = 10'b1010110000;
    16'b0000110010101100: out_v[133] = 10'b0111100011;
    16'b0010110000111000: out_v[133] = 10'b0111011110;
    16'b1000110001111100: out_v[133] = 10'b1111100001;
    16'b1000010000100100: out_v[133] = 10'b0111011110;
    16'b1000010001100100: out_v[133] = 10'b0101110001;
    16'b0000010000001100: out_v[133] = 10'b0111001001;
    16'b0000110010111100: out_v[133] = 10'b1110111111;
    16'b0000100100110000: out_v[133] = 10'b1011100111;
    16'b1010110000101100: out_v[133] = 10'b0001111110;
    16'b0100001001000000: out_v[133] = 10'b0010011111;
    16'b0000001001100000: out_v[133] = 10'b0100101011;
    16'b0110001001100000: out_v[133] = 10'b1011001011;
    16'b0000001000000000: out_v[133] = 10'b0000000110;
    16'b0000001001000000: out_v[133] = 10'b1100110001;
    16'b0000001001100100: out_v[133] = 10'b0000010111;
    16'b0100001000000000: out_v[133] = 10'b1000100111;
    16'b0010001001000000: out_v[133] = 10'b1011010111;
    16'b0010001001100100: out_v[133] = 10'b1001000101;
    16'b0000000001100000: out_v[133] = 10'b0111000010;
    16'b0010001001100000: out_v[133] = 10'b0011110011;
    16'b0100001001100000: out_v[133] = 10'b0001111001;
    16'b0000001001101100: out_v[133] = 10'b0111010111;
    16'b0100001011000000: out_v[133] = 10'b1111111111;
    16'b0010001001101100: out_v[133] = 10'b0001001111;
    16'b1100001001000000: out_v[133] = 10'b1101010010;
    16'b0100001010000000: out_v[133] = 10'b1000100010;
    16'b0010001001000100: out_v[133] = 10'b0111000101;
    16'b0100001001100100: out_v[133] = 10'b0000111001;
    16'b0010001001001100: out_v[133] = 10'b0011000101;
    16'b1000000001100000: out_v[133] = 10'b0001010110;
    16'b0100001000100000: out_v[133] = 10'b1011100101;
    16'b1100001001100000: out_v[133] = 10'b0010111011;
    16'b0100001001001100: out_v[133] = 10'b0110001101;
    16'b1000000001000000: out_v[133] = 10'b0110101101;
    16'b1100001101000000: out_v[133] = 10'b1100101111;
    16'b1100001001001000: out_v[133] = 10'b0001110111;
    16'b1100011001001100: out_v[133] = 10'b1001011100;
    16'b1000001001000001: out_v[133] = 10'b1111100111;
    16'b1100001001000001: out_v[133] = 10'b0001001001;
    16'b1000001001000000: out_v[133] = 10'b0111100001;
    16'b0110001100100001: out_v[133] = 10'b0001110111;
    16'b1100001001010000: out_v[133] = 10'b1101001101;
    16'b0100001101100000: out_v[133] = 10'b1011110000;
    16'b1100001101010000: out_v[133] = 10'b0100101001;
    16'b0100001100100000: out_v[133] = 10'b1110010110;
    16'b1100001101100000: out_v[133] = 10'b0110100101;
    16'b0100001001000001: out_v[133] = 10'b1011101001;
    16'b1100001001001100: out_v[133] = 10'b0101101010;
    16'b0000000001000000: out_v[133] = 10'b0111101010;
    16'b1100001000100000: out_v[133] = 10'b0001110000;
    16'b1000001001100000: out_v[133] = 10'b1111100000;
    16'b1100001101000001: out_v[133] = 10'b1101100111;
    16'b1100001101100001: out_v[133] = 10'b1101111010;
    16'b0100001101000000: out_v[133] = 10'b1000010111;
    16'b1100001011000000: out_v[133] = 10'b1001100011;
    16'b0100001000100001: out_v[133] = 10'b1110010001;
    16'b0100001100100001: out_v[133] = 10'b1111011011;
    16'b1010000100000000: out_v[133] = 10'b1001111000;
    16'b0000000000100000: out_v[133] = 10'b0000011101;
    16'b1010000000000000: out_v[133] = 10'b0001011000;
    16'b1000000000101100: out_v[133] = 10'b0100100011;
    16'b0010001100000000: out_v[133] = 10'b0011111001;
    16'b0110001100000000: out_v[133] = 10'b0001111110;
    16'b1000010000000000: out_v[133] = 10'b1011011111;
    16'b1000000100100000: out_v[133] = 10'b1110010011;
    16'b1010000100000001: out_v[133] = 10'b0011001111;
    16'b0000000000000000: out_v[133] = 10'b0010101001;
    16'b0010000000000000: out_v[133] = 10'b1111001011;
    16'b0010000100000000: out_v[133] = 10'b0010111100;
    16'b1000000000000000: out_v[133] = 10'b0011011110;
    16'b1010010000000000: out_v[133] = 10'b1101000101;
    16'b1000010001100000: out_v[133] = 10'b1100011111;
    16'b1000000100000000: out_v[133] = 10'b0001011111;
    16'b1010000000100000: out_v[133] = 10'b0010011011;
    16'b1010000100100000: out_v[133] = 10'b1011011011;
    16'b1000001000100000: out_v[133] = 10'b0011110111;
    16'b1010010000100000: out_v[133] = 10'b0011101011;
    16'b0000001000100000: out_v[133] = 10'b0110001000;
    16'b0000010000100000: out_v[133] = 10'b1000001110;
    16'b1000000000101000: out_v[133] = 10'b0100011111;
    16'b0010001000000000: out_v[133] = 10'b1011001011;
    16'b1010010100000000: out_v[133] = 10'b1011110111;
    16'b1110001100000000: out_v[133] = 10'b0010001011;
    16'b1000010100100000: out_v[133] = 10'b1011011011;
    16'b1110111001001000: out_v[133] = 10'b0111011100;
    16'b1110111000000000: out_v[133] = 10'b0011100111;
    16'b1100011001101100: out_v[133] = 10'b1100001110;
    16'b1010100000000000: out_v[133] = 10'b1010110111;
    16'b1100111001100000: out_v[133] = 10'b0111001011;
    16'b1110011000001100: out_v[133] = 10'b1011100110;
    16'b1000011001101100: out_v[133] = 10'b0111011011;
    16'b1110111000001000: out_v[133] = 10'b0111010111;
    16'b1110101000000000: out_v[133] = 10'b0111110011;
    16'b1100111011101000: out_v[133] = 10'b1111101111;
    16'b1100111001001100: out_v[133] = 10'b1011011110;
    16'b1100011011001100: out_v[133] = 10'b1111001010;
    16'b1110011000001000: out_v[133] = 10'b0010110001;
    16'b1110101100000000: out_v[133] = 10'b0101110111;
    16'b1100111001101100: out_v[133] = 10'b1101011111;
    16'b1110011000000000: out_v[133] = 10'b1111000011;
    16'b1100011000001100: out_v[133] = 10'b1101001010;
    16'b1100101100000001: out_v[133] = 10'b0011100101;
    16'b1100011001000000: out_v[133] = 10'b1101010100;
    16'b1100011001100000: out_v[133] = 10'b1010000011;
    16'b1100011011101100: out_v[133] = 10'b0101010011;
    16'b1000011001001100: out_v[133] = 10'b0011111111;
    16'b1100011001101000: out_v[133] = 10'b0011111011;
    16'b1100111011101100: out_v[133] = 10'b1010010111;
    16'b1100101001100000: out_v[133] = 10'b0101011011;
    16'b1000010001101000: out_v[133] = 10'b1000110111;
    16'b1100111001101000: out_v[133] = 10'b0011101011;
    16'b1100011001001000: out_v[133] = 10'b1101111011;
    16'b1000111001001100: out_v[133] = 10'b0111111111;
    16'b1110111000001100: out_v[133] = 10'b1000101010;
    16'b1110011001001100: out_v[133] = 10'b1100001100;
    16'b1110111100000000: out_v[133] = 10'b0111001100;
    16'b1010110000001000: out_v[133] = 10'b0101110010;
    16'b0100011001101100: out_v[133] = 10'b1101111000;
    16'b0000010001001100: out_v[133] = 10'b0111100011;
    16'b1010010000001000: out_v[133] = 10'b0000110101;
    16'b0000011000101100: out_v[133] = 10'b0001111110;
    16'b1000110010101100: out_v[133] = 10'b0011001110;
    16'b0000010010101100: out_v[133] = 10'b0111000111;
    16'b1000010010101100: out_v[133] = 10'b1010110110;
    16'b0000011001101100: out_v[133] = 10'b0001111010;
    16'b0110011001001100: out_v[133] = 10'b0100001101;
    16'b0000010001101100: out_v[133] = 10'b0111000000;
    16'b0100011011101100: out_v[133] = 10'b1111101011;
    16'b0000011001000000: out_v[133] = 10'b0010011011;
    16'b1000010000101000: out_v[133] = 10'b0101010111;
    16'b0100111001101100: out_v[133] = 10'b1000010111;
    16'b0000010001000000: out_v[133] = 10'b1111000110;
    16'b0100011001000000: out_v[133] = 10'b1110000100;
    16'b1100011000101100: out_v[133] = 10'b1010001110;
    16'b1000011001111100: out_v[133] = 10'b1010111001;
    16'b0100011000101100: out_v[133] = 10'b0001100110;
    16'b1100011001111100: out_v[133] = 10'b1011100110;
    16'b1100111001111100: out_v[133] = 10'b0011100011;
    16'b1100011000111100: out_v[133] = 10'b0110111110;
    16'b1000011000101100: out_v[133] = 10'b1001001111;
    16'b1000011001100100: out_v[133] = 10'b0010110101;
    16'b1100001001100100: out_v[133] = 10'b1001000110;
    16'b1000111001111100: out_v[133] = 10'b1100111110;
    16'b1100001000100100: out_v[133] = 10'b1011111001;
    16'b1100011001100100: out_v[133] = 10'b0111110111;
    16'b1100011000100100: out_v[133] = 10'b1010110111;
    16'b1000010001001100: out_v[133] = 10'b1101001111;
    16'b1000011001101000: out_v[133] = 10'b1101000010;
    16'b1000111001101100: out_v[133] = 10'b0110100101;
    16'b1000001001001100: out_v[133] = 10'b0100000111;
    16'b1000010101101100: out_v[133] = 10'b1010000011;
    16'b1000000101101100: out_v[133] = 10'b1101000011;
    16'b1010100000001100: out_v[133] = 10'b0110101111;
    16'b1000000001101100: out_v[133] = 10'b1000111110;
    16'b0000000001101100: out_v[133] = 10'b1101010101;
    16'b1000110001001100: out_v[133] = 10'b0111010010;
    16'b1010110001101100: out_v[133] = 10'b0101101101;
    16'b0000001001001100: out_v[133] = 10'b0111011100;
    16'b1000001001101100: out_v[133] = 10'b1100011001;
    16'b1000000001001100: out_v[133] = 10'b0110111110;
    16'b1010000000001100: out_v[133] = 10'b1101000010;
    16'b1000001101101100: out_v[133] = 10'b1101010101;
    16'b1100001001101100: out_v[133] = 10'b0011100110;
    16'b1000000101100000: out_v[133] = 10'b0111110101;
    16'b1010110000001100: out_v[133] = 10'b0011001110;
    16'b1000000001101000: out_v[133] = 10'b0101011011;
    16'b1000110000001100: out_v[133] = 10'b0111110010;
    16'b0000011001001100: out_v[133] = 10'b1011001101;
    16'b1000001101001100: out_v[133] = 10'b0001110111;
    16'b0100011000001100: out_v[133] = 10'b1101100110;
    16'b0110011000001100: out_v[133] = 10'b0110110110;
    16'b0100011001101000: out_v[133] = 10'b1000110011;
    16'b0100011001001100: out_v[133] = 10'b1000111100;
    16'b0100001000101100: out_v[133] = 10'b0111000000;
    16'b0100011000001000: out_v[133] = 10'b1111100110;
    16'b0110011000000000: out_v[133] = 10'b1111000011;
    16'b0110011000001000: out_v[133] = 10'b0011010111;
    16'b0100001000001100: out_v[133] = 10'b1111010001;
    16'b0100001001101100: out_v[133] = 10'b0111111011;
    16'b0100011001001000: out_v[133] = 10'b0011011001;
    16'b1110011001101100: out_v[133] = 10'b1111010011;
    16'b0100011000101000: out_v[133] = 10'b0111110111;
    16'b0110011001001000: out_v[133] = 10'b0101101011;
    16'b0110011001101100: out_v[133] = 10'b0111111110;
    16'b1110101000001000: out_v[133] = 10'b1101000111;
    16'b1110111001001100: out_v[133] = 10'b1000011101;
    16'b1000110001101000: out_v[133] = 10'b1101100001;
    16'b0000010001101000: out_v[133] = 10'b1101001100;
    16'b1100111000101100: out_v[133] = 10'b1100011000;
    16'b1110111001101100: out_v[133] = 10'b1001011111;
    default: out_v[133] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000100000000110: out_v[134] = 10'b0011011001;
    16'b0000100001010110: out_v[134] = 10'b0110010001;
    16'b0000100001000100: out_v[134] = 10'b1110110011;
    16'b0001100001000111: out_v[134] = 10'b0000100001;
    16'b0101000001010111: out_v[134] = 10'b1100011011;
    16'b0000100001010100: out_v[134] = 10'b0011010111;
    16'b0000100001000111: out_v[134] = 10'b1011000010;
    16'b0001100001010110: out_v[134] = 10'b0000110111;
    16'b0010100001010110: out_v[134] = 10'b0111001011;
    16'b0000100000010110: out_v[134] = 10'b1011010011;
    16'b0000100001000110: out_v[134] = 10'b0011011010;
    16'b0000100001010111: out_v[134] = 10'b0101001100;
    16'b0001100001110110: out_v[134] = 10'b1101110011;
    16'b0001100000000110: out_v[134] = 10'b0101001001;
    16'b0000100000110110: out_v[134] = 10'b1010110111;
    16'b0101000001000111: out_v[134] = 10'b1001100111;
    16'b0001100001000110: out_v[134] = 10'b0110000001;
    16'b0101000001010110: out_v[134] = 10'b0010111001;
    16'b0101100001010110: out_v[134] = 10'b1100010100;
    16'b0010100100110110: out_v[134] = 10'b1011001101;
    16'b0101100001010111: out_v[134] = 10'b0101011110;
    16'b0000100000000010: out_v[134] = 10'b0001111111;
    16'b0000000000000110: out_v[134] = 10'b0010010011;
    16'b0000000000110110: out_v[134] = 10'b1001001011;
    16'b0010000100110110: out_v[134] = 10'b0111011011;
    16'b0010100000110110: out_v[134] = 10'b1000110100;
    16'b0101100001000111: out_v[134] = 10'b1001100110;
    16'b0000100000000100: out_v[134] = 10'b1001110101;
    16'b0000100000010100: out_v[134] = 10'b1111011100;
    16'b0000000001000111: out_v[134] = 10'b1011100001;
    16'b0101000000000111: out_v[134] = 10'b1010100101;
    16'b0100000000000010: out_v[134] = 10'b0001100110;
    16'b0101000000000000: out_v[134] = 10'b1101110000;
    16'b0101000001000110: out_v[134] = 10'b0101110100;
    16'b0101000000000110: out_v[134] = 10'b0010100011;
    16'b0101000000000010: out_v[134] = 10'b1011000100;
    16'b0100000001000000: out_v[134] = 10'b1100010111;
    16'b0100100001000000: out_v[134] = 10'b1011100111;
    16'b0000000001000000: out_v[134] = 10'b1010010011;
    16'b0101000000000100: out_v[134] = 10'b1011111000;
    16'b0000100001000000: out_v[134] = 10'b1010101011;
    16'b0000000000000000: out_v[134] = 10'b1100001110;
    16'b0101000000000001: out_v[134] = 10'b0010011001;
    16'b0100000000000000: out_v[134] = 10'b1101011111;
    16'b0101000000000101: out_v[134] = 10'b0110110110;
    16'b0001000000000000: out_v[134] = 10'b1001111011;
    16'b0100000000000110: out_v[134] = 10'b1110110000;
    16'b0101100001000000: out_v[134] = 10'b1001111010;
    16'b0101000001000000: out_v[134] = 10'b0000101111;
    16'b0101000001000010: out_v[134] = 10'b1100110000;
    16'b0101100001000010: out_v[134] = 10'b1100110100;
    16'b0101100001000110: out_v[134] = 10'b0111100100;
    16'b0100000001000010: out_v[134] = 10'b0111001101;
    16'b0101100000000111: out_v[134] = 10'b0111011100;
    16'b0101100001100110: out_v[134] = 10'b0110100100;
    16'b0101100001000101: out_v[134] = 10'b0110001111;
    16'b0101000000000011: out_v[134] = 10'b0110001000;
    16'b0111100001000111: out_v[134] = 10'b0101011000;
    16'b0101100001010101: out_v[134] = 10'b0111111011;
    16'b0101000000010111: out_v[134] = 10'b1101100101;
    16'b0111100101100111: out_v[134] = 10'b1110100001;
    16'b0101100001000001: out_v[134] = 10'b0000010111;
    16'b0101100001100111: out_v[134] = 10'b1011110000;
    16'b0101000001000101: out_v[134] = 10'b1001011000;
    16'b0111100101000111: out_v[134] = 10'b0000101110;
    16'b1101100001000111: out_v[134] = 10'b1111011000;
    16'b0111100101100110: out_v[134] = 10'b0111101011;
    16'b1101100001000110: out_v[134] = 10'b0111101011;
    16'b0101000000100111: out_v[134] = 10'b1010010111;
    16'b0111100100000111: out_v[134] = 10'b1101010000;
    16'b1101100001100111: out_v[134] = 10'b1110111010;
    16'b0101000001100111: out_v[134] = 10'b1001001011;
    16'b0111000100000111: out_v[134] = 10'b1001111111;
    16'b0101100001100101: out_v[134] = 10'b1010101011;
    16'b0101100001000100: out_v[134] = 10'b1011001000;
    16'b0010100100000111: out_v[134] = 10'b0011111011;
    16'b0000100001000010: out_v[134] = 10'b1001101100;
    16'b0010100101000111: out_v[134] = 10'b0011111011;
    16'b0000000000000111: out_v[134] = 10'b1101000000;
    16'b0000100000000011: out_v[134] = 10'b1101110001;
    16'b0000100000000111: out_v[134] = 10'b0101111001;
    16'b0010100100000011: out_v[134] = 10'b1101101011;
    16'b0000100001000101: out_v[134] = 10'b0100000111;
    16'b0010000100000011: out_v[134] = 10'b1011101101;
    16'b0000000001000110: out_v[134] = 10'b1101101100;
    16'b0010000100000111: out_v[134] = 10'b1000001101;
    16'b0010100100100111: out_v[134] = 10'b0111110000;
    16'b0010100000000111: out_v[134] = 10'b0111010100;
    16'b0010100001000111: out_v[134] = 10'b1010100110;
    16'b0000100001000001: out_v[134] = 10'b0110111111;
    16'b0000100000000101: out_v[134] = 10'b0100011001;
    16'b0010000100100111: out_v[134] = 10'b0100101010;
    16'b0010100101000110: out_v[134] = 10'b1101111011;
    16'b0000100000000001: out_v[134] = 10'b0110110011;
    16'b0000100001000011: out_v[134] = 10'b0101000011;
    16'b0100100001000110: out_v[134] = 10'b0011111010;
    16'b0000000001000001: out_v[134] = 10'b0110011000;
    16'b0101000001010001: out_v[134] = 10'b0100110011;
    16'b0101000001000001: out_v[134] = 10'b0111100001;
    16'b0100000001000001: out_v[134] = 10'b0001011101;
    16'b0000000000000001: out_v[134] = 10'b0100100111;
    16'b0101000000010001: out_v[134] = 10'b1010001111;
    16'b0100000000000101: out_v[134] = 10'b0010111001;
    16'b0010100001000001: out_v[134] = 10'b0101001101;
    16'b0100000001000111: out_v[134] = 10'b1100000100;
    16'b0000000001010001: out_v[134] = 10'b1111001011;
    16'b0100100001000111: out_v[134] = 10'b1000110110;
    16'b0000000001000101: out_v[134] = 10'b1011100001;
    16'b0000100001010001: out_v[134] = 10'b1001111010;
    16'b0100000000000001: out_v[134] = 10'b0000010101;
    16'b0100100001000001: out_v[134] = 10'b0110010000;
    16'b0010100101000001: out_v[134] = 10'b1110100010;
    16'b0100000001000101: out_v[134] = 10'b0001011110;
    16'b0101100001010001: out_v[134] = 10'b0101110000;
    16'b0100100001010001: out_v[134] = 10'b0101111010;
    16'b0100000001010001: out_v[134] = 10'b0101100011;
    16'b0100100001000101: out_v[134] = 10'b0110110011;
    16'b0101000000010000: out_v[134] = 10'b1000111001;
    16'b0101000001010000: out_v[134] = 10'b1011111011;
    16'b0100000001000110: out_v[134] = 10'b0011100111;
    16'b0101100011000001: out_v[134] = 10'b1000111100;
    16'b1101100001000000: out_v[134] = 10'b1011101100;
    16'b1101100001000001: out_v[134] = 10'b1011100011;
    16'b0101100011000000: out_v[134] = 10'b1001001011;
    16'b0101100000000001: out_v[134] = 10'b1010011101;
    16'b0001100001000001: out_v[134] = 10'b1101101000;
    16'b0101100011100001: out_v[134] = 10'b1110111111;
    16'b0001100011000001: out_v[134] = 10'b1010101001;
    16'b1101100001100001: out_v[134] = 10'b0111001011;
    16'b0101100011000111: out_v[134] = 10'b0111010101;
    16'b0001100000000001: out_v[134] = 10'b1111010110;
    16'b0001100001000101: out_v[134] = 10'b1111110100;
    16'b0001100001000000: out_v[134] = 10'b1101000110;
    16'b0101000011000001: out_v[134] = 10'b1110101011;
    16'b1101100001010001: out_v[134] = 10'b1111100010;
    16'b0111000101010011: out_v[134] = 10'b1001111001;
    16'b0101000001000011: out_v[134] = 10'b1001110000;
    16'b0110100101000001: out_v[134] = 10'b1111100111;
    16'b0010000001000011: out_v[134] = 10'b0001110111;
    16'b0010100101000011: out_v[134] = 10'b0111010111;
    16'b0000000001000011: out_v[134] = 10'b1001000110;
    16'b0111000000000011: out_v[134] = 10'b1101100111;
    16'b0100000000000011: out_v[134] = 10'b1101101001;
    16'b0110000101000001: out_v[134] = 10'b0111100110;
    16'b0010100100000000: out_v[134] = 10'b0111010111;
    16'b0111000001000011: out_v[134] = 10'b1111011011;
    16'b0101000001010011: out_v[134] = 10'b0100011001;
    16'b0111000101000111: out_v[134] = 10'b1011100010;
    16'b0111000100000011: out_v[134] = 10'b0010111111;
    16'b0010000101000011: out_v[134] = 10'b0110100010;
    16'b0100000001000011: out_v[134] = 10'b1011011101;
    16'b0010100101000000: out_v[134] = 10'b1010011001;
    16'b0110000101000011: out_v[134] = 10'b1101111011;
    16'b0111000101000011: out_v[134] = 10'b0101011111;
    16'b0010000101000001: out_v[134] = 10'b0111101101;
    16'b0010100101010001: out_v[134] = 10'b0001111110;
    16'b0101000000010011: out_v[134] = 10'b0110001011;
    16'b0110100101000011: out_v[134] = 10'b0011110011;
    16'b0000100001010000: out_v[134] = 10'b0110001111;
    16'b0010100001000011: out_v[134] = 10'b1000001111;
    16'b0111100001010111: out_v[134] = 10'b1011100110;
    16'b0000000001010111: out_v[134] = 10'b1101000111;
    16'b0100000001010111: out_v[134] = 10'b1011001111;
    16'b0101100000000110: out_v[134] = 10'b1101000111;
    16'b0100100001010111: out_v[134] = 10'b1111101010;
    16'b0101000000010110: out_v[134] = 10'b0100001010;
    16'b0100000000010111: out_v[134] = 10'b1000101111;
    16'b0111100101010111: out_v[134] = 10'b0100000111;
    16'b0100000000000111: out_v[134] = 10'b0001011000;
    16'b0101100001000011: out_v[134] = 10'b1100011011;
    16'b0100100001000011: out_v[134] = 10'b1001111011;
    16'b0000000000000011: out_v[134] = 10'b1111110111;
    default: out_v[134] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0110110010100000: out_v[135] = 10'b0001100100;
    16'b1011010010110000: out_v[135] = 10'b1000001111;
    16'b0100100000000000: out_v[135] = 10'b1111000001;
    16'b1001000010010000: out_v[135] = 10'b1111011101;
    16'b1001000000010000: out_v[135] = 10'b0011010001;
    16'b1101000010010000: out_v[135] = 10'b0000011111;
    16'b0000100010100000: out_v[135] = 10'b0110111011;
    16'b1101100010000000: out_v[135] = 10'b0011111101;
    16'b1101001000010000: out_v[135] = 10'b0001100001;
    16'b0100100010000000: out_v[135] = 10'b1001011010;
    16'b1101100010010000: out_v[135] = 10'b1000101111;
    16'b1101100000000000: out_v[135] = 10'b0010010101;
    16'b1111110010110000: out_v[135] = 10'b1110100101;
    16'b0000110010000000: out_v[135] = 10'b1001100001;
    16'b0000110010100000: out_v[135] = 10'b1001010101;
    16'b1011000010100000: out_v[135] = 10'b1010100011;
    16'b0010010010100000: out_v[135] = 10'b0101011100;
    16'b0010100010100000: out_v[135] = 10'b1100101010;
    16'b1111000010010000: out_v[135] = 10'b1000100011;
    16'b1101000000010000: out_v[135] = 10'b1010100011;
    16'b1111000010100000: out_v[135] = 10'b1111000010;
    16'b1111000010110000: out_v[135] = 10'b1100001011;
    16'b0000100000000000: out_v[135] = 10'b0001111001;
    16'b1011000010110000: out_v[135] = 10'b0010010000;
    16'b1011000010010000: out_v[135] = 10'b0011100000;
    16'b1111010010110000: out_v[135] = 10'b1111000011;
    16'b0000100010000000: out_v[135] = 10'b0111001101;
    16'b1101100000010000: out_v[135] = 10'b0100111110;
    16'b1101001010010000: out_v[135] = 10'b1010111110;
    16'b0010110010100000: out_v[135] = 10'b1001001111;
    16'b1101000010000000: out_v[135] = 10'b0111001011;
    16'b1001100010010000: out_v[135] = 10'b0111010011;
    16'b1011000010110100: out_v[135] = 10'b0111011001;
    16'b1101001000000000: out_v[135] = 10'b0000011011;
    16'b1100100000000000: out_v[135] = 10'b1100000011;
    16'b1001001000010000: out_v[135] = 10'b1111110101;
    16'b1101101000000000: out_v[135] = 10'b0111100101;
    16'b0100110010000000: out_v[135] = 10'b0111011001;
    16'b1001100000010000: out_v[135] = 10'b1100101110;
    16'b1111011010110000: out_v[135] = 10'b1000111111;
    16'b0010000010100000: out_v[135] = 10'b1010100010;
    16'b1101101010000000: out_v[135] = 10'b1111000110;
    16'b1011100010110000: out_v[135] = 10'b0010011001;
    16'b1111100010110000: out_v[135] = 10'b0001011111;
    16'b1101101000010000: out_v[135] = 10'b1110111110;
    16'b1111001010110000: out_v[135] = 10'b1111001111;
    16'b1101101010010000: out_v[135] = 10'b1011011110;
    16'b0100110010100000: out_v[135] = 10'b0111110010;
    16'b0110100010100000: out_v[135] = 10'b0101001000;
    16'b1111100010100000: out_v[135] = 10'b1011000110;
    16'b0100000000000000: out_v[135] = 10'b0110000010;
    16'b0000000000000000: out_v[135] = 10'b1101001110;
    16'b0000010000000000: out_v[135] = 10'b0010110010;
    16'b0000000010100000: out_v[135] = 10'b1110000001;
    16'b0000000010000000: out_v[135] = 10'b1100000111;
    16'b0100010000000000: out_v[135] = 10'b0101001100;
    16'b0000010010100000: out_v[135] = 10'b0100111001;
    16'b0010000010000000: out_v[135] = 10'b0000100110;
    16'b0010000010000100: out_v[135] = 10'b1000100110;
    16'b1001100000000000: out_v[135] = 10'b0011101110;
    16'b0000000000000100: out_v[135] = 10'b0100100100;
    16'b0110000010100000: out_v[135] = 10'b0001110110;
    16'b0110000000000000: out_v[135] = 10'b0011110010;
    16'b0000000000010000: out_v[135] = 10'b0000110101;
    16'b1001100000000100: out_v[135] = 10'b0100000111;
    16'b1001000000000100: out_v[135] = 10'b1001001100;
    16'b0110000010000000: out_v[135] = 10'b0001010111;
    16'b0010000000000000: out_v[135] = 10'b1010000110;
    16'b0000100000000100: out_v[135] = 10'b0010100100;
    16'b1101100000000100: out_v[135] = 10'b1111101001;
    16'b0000001000000000: out_v[135] = 10'b0000101010;
    16'b0100000001000000: out_v[135] = 10'b1000011101;
    16'b1001000000000000: out_v[135] = 10'b1001101100;
    16'b1001001000000000: out_v[135] = 10'b1100001111;
    16'b0100000000000100: out_v[135] = 10'b1111011111;
    16'b1111101000000000: out_v[135] = 10'b0000110110;
    16'b0100000010000000: out_v[135] = 10'b0101010011;
    16'b0010100010000000: out_v[135] = 10'b0001011001;
    16'b0110010010100000: out_v[135] = 10'b1010110110;
    16'b1001101000000000: out_v[135] = 10'b1011000111;
    16'b0010100000000000: out_v[135] = 10'b1011010011;
    16'b0010000010100100: out_v[135] = 10'b0010111110;
    16'b0100001000000000: out_v[135] = 10'b0100011000;
    16'b0000100000010000: out_v[135] = 10'b1001001110;
    16'b0100100011000000: out_v[135] = 10'b0011111110;
    16'b0100100001000000: out_v[135] = 10'b0110001000;
    16'b0100101010000000: out_v[135] = 10'b1001011011;
    16'b0100010010000000: out_v[135] = 10'b1011011100;
    16'b0000010010000000: out_v[135] = 10'b1011001011;
    16'b0100010010100000: out_v[135] = 10'b0111101011;
    16'b0100001010000000: out_v[135] = 10'b0111110100;
    16'b0110110011100000: out_v[135] = 10'b0110010110;
    16'b0100101000000000: out_v[135] = 10'b0010111100;
    16'b0000110000000000: out_v[135] = 10'b1010010011;
    16'b1011000000000000: out_v[135] = 10'b0010111000;
    16'b0100110000000000: out_v[135] = 10'b1001011110;
    16'b1011100010100000: out_v[135] = 10'b0111111011;
    16'b1001110000000000: out_v[135] = 10'b0101111011;
    16'b0100100010100000: out_v[135] = 10'b0001011111;
    16'b1101100010100000: out_v[135] = 10'b0100111001;
    16'b1000100000000000: out_v[135] = 10'b0110011100;
    16'b1001100010100000: out_v[135] = 10'b0110010000;
    16'b1101000000000000: out_v[135] = 10'b1000111011;
    16'b1101110000000000: out_v[135] = 10'b1111001010;
    16'b1011100000000000: out_v[135] = 10'b0000111011;
    16'b1001110010100000: out_v[135] = 10'b0011100100;
    16'b1001000010100000: out_v[135] = 10'b1100010101;
    16'b0110100010000000: out_v[135] = 10'b0100101001;
    16'b0000100100000000: out_v[135] = 10'b0011110100;
    16'b1111110010100000: out_v[135] = 10'b1010111000;
    16'b0000101000000000: out_v[135] = 10'b0010101000;
    16'b1000000000010000: out_v[135] = 10'b1011111110;
    16'b0010100010010000: out_v[135] = 10'b0001001010;
    16'b0000100010010000: out_v[135] = 10'b1100101011;
    16'b1000100000010000: out_v[135] = 10'b1001010111;
    16'b0010010000100000: out_v[135] = 10'b0101001001;
    16'b0010110000100000: out_v[135] = 10'b0110000011;
    16'b0100000010100000: out_v[135] = 10'b0010111101;
    default: out_v[135] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1000000000010000: out_v[136] = 10'b1101001101;
    16'b1000011010000000: out_v[136] = 10'b0000011010;
    16'b0001011010000000: out_v[136] = 10'b1111011011;
    16'b1000001010000000: out_v[136] = 10'b0001111001;
    16'b0000001000010000: out_v[136] = 10'b1110110001;
    16'b1000001010000010: out_v[136] = 10'b1011101010;
    16'b0000011010000010: out_v[136] = 10'b1001111010;
    16'b0000000010000000: out_v[136] = 10'b1101101011;
    16'b0000011010000000: out_v[136] = 10'b0111000111;
    16'b1000001000010000: out_v[136] = 10'b1001101101;
    16'b1000011010010000: out_v[136] = 10'b0110010101;
    16'b0000001010000010: out_v[136] = 10'b0010110001;
    16'b1000001010010010: out_v[136] = 10'b0010111101;
    16'b1000011010000010: out_v[136] = 10'b0000111011;
    16'b1000010010000000: out_v[136] = 10'b1011110011;
    16'b1000001010010000: out_v[136] = 10'b1111010100;
    16'b0000001010010000: out_v[136] = 10'b0101000110;
    16'b1001001010010010: out_v[136] = 10'b0110101001;
    16'b0000000010000010: out_v[136] = 10'b1001110111;
    16'b1001001010000000: out_v[136] = 10'b1011011100;
    16'b1001011010000000: out_v[136] = 10'b0100001010;
    16'b1000000010000000: out_v[136] = 10'b0101100101;
    16'b0000010010010010: out_v[136] = 10'b0110001011;
    16'b1000011010010010: out_v[136] = 10'b0000110111;
    16'b0000001010000000: out_v[136] = 10'b1110000101;
    16'b1000001000010010: out_v[136] = 10'b1001100111;
    16'b1001001010000010: out_v[136] = 10'b1011011000;
    16'b0001001010000000: out_v[136] = 10'b0011100110;
    16'b0000010010000010: out_v[136] = 10'b1100100111;
    16'b0000001000010010: out_v[136] = 10'b1001001110;
    16'b0000000000010000: out_v[136] = 10'b0100011111;
    16'b1000001000000000: out_v[136] = 10'b1000101010;
    16'b0000001000000000: out_v[136] = 10'b0000111010;
    16'b0000011010010010: out_v[136] = 10'b1010011110;
    16'b1000011000000000: out_v[136] = 10'b0111010010;
    16'b1001011010000010: out_v[136] = 10'b0111011111;
    16'b1000010010000010: out_v[136] = 10'b0100001011;
    16'b0000001010010010: out_v[136] = 10'b0010001110;
    16'b0000000000010010: out_v[136] = 10'b0010011101;
    16'b0000000000000010: out_v[136] = 10'b0111110000;
    16'b1000001000000010: out_v[136] = 10'b0110001111;
    16'b0000001000000010: out_v[136] = 10'b0110100111;
    16'b1000000000000010: out_v[136] = 10'b0111000000;
    16'b0000000000000000: out_v[136] = 10'b0010010000;
    16'b0000000010010010: out_v[136] = 10'b1100100111;
    16'b1000000000000000: out_v[136] = 10'b1001101101;
    16'b1000000000010010: out_v[136] = 10'b1000011110;
    16'b1000000010010010: out_v[136] = 10'b0010010101;
    16'b1001001000000011: out_v[136] = 10'b0100011111;
    16'b1000000010000010: out_v[136] = 10'b1001001110;
    16'b1001001000010010: out_v[136] = 10'b0010100011;
    16'b1001000010010010: out_v[136] = 10'b0000011110;
    16'b0001001000010000: out_v[136] = 10'b0010011110;
    16'b1001001010010011: out_v[136] = 10'b1000100111;
    16'b1000000010010011: out_v[136] = 10'b0111001111;
    16'b0001000010010010: out_v[136] = 10'b0000110111;
    16'b0001001000000010: out_v[136] = 10'b0110000101;
    16'b1001001000000010: out_v[136] = 10'b1100110110;
    16'b0001001000010010: out_v[136] = 10'b0111000010;
    16'b0001001010010010: out_v[136] = 10'b1111001011;
    16'b0001000000010010: out_v[136] = 10'b1101100101;
    16'b1001001000010011: out_v[136] = 10'b1111010001;
    16'b1000010010010010: out_v[136] = 10'b0101100110;
    16'b0000000010010000: out_v[136] = 10'b0000010110;
    16'b0000000010011010: out_v[136] = 10'b1111100101;
    16'b0001001010010000: out_v[136] = 10'b1010011111;
    16'b0000000010010011: out_v[136] = 10'b0110010000;
    16'b1001000000010010: out_v[136] = 10'b0010111010;
    16'b1000000010010000: out_v[136] = 10'b0100010011;
    16'b1001000000000000: out_v[136] = 10'b1001001100;
    16'b1000000000000001: out_v[136] = 10'b0001011001;
    16'b1001001000010000: out_v[136] = 10'b1011110111;
    16'b0001000000000000: out_v[136] = 10'b1010011000;
    16'b0001001000000000: out_v[136] = 10'b0100010010;
    16'b1001000000000001: out_v[136] = 10'b0010111010;
    16'b1001001000000001: out_v[136] = 10'b0001110110;
    16'b1001001000000000: out_v[136] = 10'b1111011010;
    16'b1001000000010000: out_v[136] = 10'b0010111011;
    16'b0000011000010000: out_v[136] = 10'b1100101111;
    16'b0000011000000000: out_v[136] = 10'b0011000100;
    16'b1000011000000010: out_v[136] = 10'b0100011111;
    16'b0000010000000010: out_v[136] = 10'b1011000011;
    16'b0001000000010001: out_v[136] = 10'b0110110000;
    16'b0001011000010000: out_v[136] = 10'b0010000111;
    16'b0000010000010010: out_v[136] = 10'b1000110000;
    16'b0000000000010001: out_v[136] = 10'b1100110101;
    16'b0000011000000010: out_v[136] = 10'b1011101111;
    16'b0000011000010010: out_v[136] = 10'b1101101001;
    16'b1000010000000010: out_v[136] = 10'b0111011110;
    16'b0001000000010000: out_v[136] = 10'b1110010011;
    16'b0001000000000001: out_v[136] = 10'b1110100011;
    16'b0000010000010000: out_v[136] = 10'b1000101011;
    16'b0000000000000001: out_v[136] = 10'b1010011010;
    16'b1000011000010010: out_v[136] = 10'b1101011000;
    16'b0000010000000000: out_v[136] = 10'b1001111010;
    16'b1000011000010000: out_v[136] = 10'b1011001110;
    16'b1000010000000000: out_v[136] = 10'b0010101011;
    16'b1000001000011010: out_v[136] = 10'b0001111010;
    16'b0000001000011010: out_v[136] = 10'b1001000001;
    16'b1000001010011010: out_v[136] = 10'b1110011011;
    16'b0000000000011010: out_v[136] = 10'b0011101110;
    16'b0000001010001010: out_v[136] = 10'b1000011011;
    16'b0001011000000010: out_v[136] = 10'b1101001011;
    16'b0000000100000000: out_v[136] = 10'b0111011110;
    16'b1001000100000000: out_v[136] = 10'b0101110101;
    16'b0001001100000000: out_v[136] = 10'b0000100111;
    16'b1001001100000000: out_v[136] = 10'b0100010100;
    16'b0000001100000000: out_v[136] = 10'b1001001010;
    16'b0001000000000010: out_v[136] = 10'b0111000000;
    16'b1001000000000010: out_v[136] = 10'b0010101100;
    16'b0001000100000000: out_v[136] = 10'b0111010010;
    16'b1001011000000010: out_v[136] = 10'b0011100111;
    16'b1000001100000000: out_v[136] = 10'b1100001000;
    16'b0001010000000010: out_v[136] = 10'b0111111011;
    16'b1000010000010000: out_v[136] = 10'b1111011001;
    16'b1000010000010010: out_v[136] = 10'b0011111000;
    16'b0000011010010000: out_v[136] = 10'b1110010010;
    16'b1000010010010000: out_v[136] = 10'b0110000101;
    16'b1001011000010010: out_v[136] = 10'b1000001100;
    16'b1000000100000000: out_v[136] = 10'b1101100111;
    16'b1000000100010000: out_v[136] = 10'b1010001011;
    16'b1000000000010001: out_v[136] = 10'b0010101111;
    16'b1000001100010000: out_v[136] = 10'b1101100101;
    16'b1001000000010001: out_v[136] = 10'b1001110111;
    16'b1001000000010011: out_v[136] = 10'b1100101010;
    default: out_v[136] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1000000000000000: out_v[137] = 10'b1001001011;
    16'b1000100110000011: out_v[137] = 10'b1011000010;
    16'b1000100010000011: out_v[137] = 10'b1110010110;
    16'b1000000100000000: out_v[137] = 10'b1011001100;
    16'b0000100000000011: out_v[137] = 10'b1001010101;
    16'b0000100010000001: out_v[137] = 10'b0001110011;
    16'b0000000000000000: out_v[137] = 10'b0010010110;
    16'b1000100010000000: out_v[137] = 10'b0110110001;
    16'b1000100110000000: out_v[137] = 10'b1111111110;
    16'b1000000101000000: out_v[137] = 10'b0101010000;
    16'b1000100010000001: out_v[137] = 10'b1100111010;
    16'b1000000010000000: out_v[137] = 10'b1010011001;
    16'b1000000010000001: out_v[137] = 10'b1000110111;
    16'b1000100000000001: out_v[137] = 10'b1001000011;
    16'b1000101010000000: out_v[137] = 10'b1111000011;
    16'b1000100000000011: out_v[137] = 10'b1000100001;
    16'b1000000110000000: out_v[137] = 10'b1001111010;
    16'b0000100010000011: out_v[137] = 10'b0000000101;
    16'b1000000000000001: out_v[137] = 10'b0111100001;
    16'b1010100010000011: out_v[137] = 10'b1010011011;
    16'b0000100000000001: out_v[137] = 10'b1111111010;
    16'b1000001111000000: out_v[137] = 10'b1000010111;
    16'b0000000101000000: out_v[137] = 10'b1010001001;
    16'b1000101010000011: out_v[137] = 10'b1101000011;
    16'b1000100110000001: out_v[137] = 10'b1011001111;
    16'b1000100100000001: out_v[137] = 10'b1101001011;
    16'b1000100111000011: out_v[137] = 10'b1000000011;
    16'b1000101111000000: out_v[137] = 10'b0000011111;
    16'b1000000111000000: out_v[137] = 10'b1010000111;
    16'b1000100111000000: out_v[137] = 10'b1010010101;
    16'b0010100010000011: out_v[137] = 10'b1011110101;
    16'b1000101111000001: out_v[137] = 10'b1010110011;
    16'b1000101110000000: out_v[137] = 10'b1110101110;
    16'b1000100111000001: out_v[137] = 10'b1001010010;
    16'b1000100000000000: out_v[137] = 10'b0011001110;
    16'b0000100010000000: out_v[137] = 10'b1101000101;
    16'b1000100101000000: out_v[137] = 10'b0100010100;
    16'b1000101010000001: out_v[137] = 10'b0001110111;
    16'b0000000000000001: out_v[137] = 10'b1110101000;
    16'b0000001000000000: out_v[137] = 10'b1101101110;
    16'b0000000100000000: out_v[137] = 10'b1100001110;
    16'b0000000100000001: out_v[137] = 10'b0000101111;
    16'b0000100100000000: out_v[137] = 10'b0100100111;
    16'b0010000101000000: out_v[137] = 10'b1000000111;
    16'b0000000101000001: out_v[137] = 10'b1001110000;
    16'b1000100111010000: out_v[137] = 10'b1011101010;
    16'b0000100101000000: out_v[137] = 10'b1011000110;
    16'b1010000101000000: out_v[137] = 10'b1110110100;
    16'b1000000101000001: out_v[137] = 10'b1010110100;
    16'b0000001111000000: out_v[137] = 10'b0101000100;
    16'b0010000100000000: out_v[137] = 10'b1100110101;
    16'b0000000111000000: out_v[137] = 10'b0010110010;
    16'b0010000000000000: out_v[137] = 10'b1000001010;
    16'b0010000101000001: out_v[137] = 10'b1001111011;
    16'b0000000001000000: out_v[137] = 10'b1111011000;
    16'b1010000000000001: out_v[137] = 10'b0100110001;
    16'b1010000000000000: out_v[137] = 10'b0010001000;
    16'b0000000010000000: out_v[137] = 10'b0001011110;
    16'b0000000001000001: out_v[137] = 10'b0110100001;
    16'b1000000000010000: out_v[137] = 10'b0111011111;
    16'b0000001101000000: out_v[137] = 10'b0010110000;
    16'b0000100101000001: out_v[137] = 10'b0011010001;
    16'b0000100111000000: out_v[137] = 10'b1010101010;
    16'b1000100101000001: out_v[137] = 10'b1001001010;
    16'b0000101111000001: out_v[137] = 10'b1111010010;
    16'b1000100101000011: out_v[137] = 10'b1001111000;
    16'b0000101101000000: out_v[137] = 10'b0101010000;
    16'b0000100001000001: out_v[137] = 10'b0111011011;
    16'b0000000111000001: out_v[137] = 10'b0111011010;
    16'b0000001100000000: out_v[137] = 10'b0101010100;
    16'b1000100001000001: out_v[137] = 10'b1111001111;
    16'b1010100000000010: out_v[137] = 10'b1101110001;
    16'b1000101101000001: out_v[137] = 10'b1010110010;
    16'b0000100101000011: out_v[137] = 10'b1101010010;
    16'b1000101111000011: out_v[137] = 10'b1011011001;
    16'b1000101101000000: out_v[137] = 10'b1111101000;
    16'b0000101111000000: out_v[137] = 10'b1011001111;
    16'b0000100111000001: out_v[137] = 10'b1110110100;
    16'b1000001000000001: out_v[137] = 10'b1001110110;
    16'b0000000110000000: out_v[137] = 10'b0100100000;
    16'b0000001000000001: out_v[137] = 10'b0011110110;
    16'b0000001101000001: out_v[137] = 10'b1110001011;
    16'b0000001001000000: out_v[137] = 10'b1100011011;
    16'b1000001000000000: out_v[137] = 10'b1000110111;
    16'b0000000010000001: out_v[137] = 10'b0110100001;
    16'b1000001100000000: out_v[137] = 10'b0010100011;
    16'b0000000110000001: out_v[137] = 10'b1111001010;
    16'b0000001001000001: out_v[137] = 10'b1111111001;
    16'b1000000100000001: out_v[137] = 10'b0111001110;
    16'b0000100100000001: out_v[137] = 10'b0011101010;
    16'b1000100100000000: out_v[137] = 10'b0011010110;
    16'b1010000111000001: out_v[137] = 10'b1111100000;
    16'b0010000000000001: out_v[137] = 10'b1001110110;
    16'b1010000101000001: out_v[137] = 10'b1011100100;
    16'b0010000100000001: out_v[137] = 10'b1000001110;
    16'b1000000111000001: out_v[137] = 10'b1111010010;
    16'b0010000111000001: out_v[137] = 10'b0011000001;
    16'b0000000101000011: out_v[137] = 10'b0000111101;
    16'b1010000111000011: out_v[137] = 10'b1010101111;
    16'b1000000111000011: out_v[137] = 10'b0111001111;
    16'b0000001010000000: out_v[137] = 10'b1011011110;
    16'b0000000011000000: out_v[137] = 10'b0111111010;
    16'b0000000011000001: out_v[137] = 10'b1110110111;
    16'b0000001111000001: out_v[137] = 10'b1111101111;
    16'b0000001110000000: out_v[137] = 10'b1011111010;
    16'b0000001110000001: out_v[137] = 10'b1111001111;
    16'b0000100111000011: out_v[137] = 10'b1000110010;
    16'b1010100101000011: out_v[137] = 10'b1010001110;
    16'b1010100000000011: out_v[137] = 10'b1011010111;
    default: out_v[137] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100000000101011: out_v[138] = 10'b0100000101;
    16'b0100010000100010: out_v[138] = 10'b1010111110;
    16'b0000000000100000: out_v[138] = 10'b1011010101;
    16'b0000100000001011: out_v[138] = 10'b1010100010;
    16'b0000010000101011: out_v[138] = 10'b0001001001;
    16'b0000100000101011: out_v[138] = 10'b0110000101;
    16'b0100010000000000: out_v[138] = 10'b1110100111;
    16'b0000010000001011: out_v[138] = 10'b0110101101;
    16'b0000010000000000: out_v[138] = 10'b1011000111;
    16'b0000100000001010: out_v[138] = 10'b1000001110;
    16'b0100000000100011: out_v[138] = 10'b0101010011;
    16'b0000000000100011: out_v[138] = 10'b0100010011;
    16'b0100000000100010: out_v[138] = 10'b1011011111;
    16'b0000000000101011: out_v[138] = 10'b0111110001;
    16'b0000000000101010: out_v[138] = 10'b1110010111;
    16'b0100000000100000: out_v[138] = 10'b0011110110;
    16'b0100010000100000: out_v[138] = 10'b1111100110;
    16'b0000000000100010: out_v[138] = 10'b1011001111;
    16'b0000010000100010: out_v[138] = 10'b1101101111;
    16'b0000010000100011: out_v[138] = 10'b0001001110;
    16'b0000010000101010: out_v[138] = 10'b1100000111;
    16'b0100010000101010: out_v[138] = 10'b0011111111;
    16'b0100010000101011: out_v[138] = 10'b0000001001;
    16'b0000010000101000: out_v[138] = 10'b0001101011;
    16'b0000000000001011: out_v[138] = 10'b0010101010;
    16'b0100010000100011: out_v[138] = 10'b0011000011;
    16'b0100100000100011: out_v[138] = 10'b1101011010;
    16'b0100100000001011: out_v[138] = 10'b1001101001;
    16'b0000000000101000: out_v[138] = 10'b0011011011;
    16'b0000010000000011: out_v[138] = 10'b0100011110;
    16'b0100100000101011: out_v[138] = 10'b1110000001;
    16'b0100010000001011: out_v[138] = 10'b1001010011;
    16'b0000010000100000: out_v[138] = 10'b0011100011;
    16'b0000010000000010: out_v[138] = 10'b1100000100;
    16'b0000100000100011: out_v[138] = 10'b0110011001;
    16'b0000000000001000: out_v[138] = 10'b0100011011;
    16'b0100000000101010: out_v[138] = 10'b0111100111;
    16'b0000100000001000: out_v[138] = 10'b0100011111;
    16'b0000000000000000: out_v[138] = 10'b0001110010;
    16'b0100000000001001: out_v[138] = 10'b1001000010;
    16'b0000000000000011: out_v[138] = 10'b0101011110;
    16'b0100000000001011: out_v[138] = 10'b0010110010;
    16'b0100000000001000: out_v[138] = 10'b1001001011;
    16'b0000000000001001: out_v[138] = 10'b1110100000;
    16'b0000000000000001: out_v[138] = 10'b1100001101;
    16'b0000100000000000: out_v[138] = 10'b0001110010;
    16'b0100000000001010: out_v[138] = 10'b0110101100;
    16'b0000000000001010: out_v[138] = 10'b1111001000;
    16'b0100100000000000: out_v[138] = 10'b0010100010;
    16'b0000100000100000: out_v[138] = 10'b1100011000;
    16'b0100100000001000: out_v[138] = 10'b1001000101;
    16'b0100100000100000: out_v[138] = 10'b0110011010;
    16'b0100100000001010: out_v[138] = 10'b1111011010;
    16'b0100000000000000: out_v[138] = 10'b0100101010;
    16'b0000100000100010: out_v[138] = 10'b1110101000;
    16'b0000100000000010: out_v[138] = 10'b1011100000;
    16'b0000000000000010: out_v[138] = 10'b0011101000;
    16'b0000100000101000: out_v[138] = 10'b0110011110;
    16'b0000110000001011: out_v[138] = 10'b0010111110;
    16'b0100100000100010: out_v[138] = 10'b1101111001;
    16'b0100100000001001: out_v[138] = 10'b1110011110;
    16'b0100000000000011: out_v[138] = 10'b1100011100;
    16'b0101100000001010: out_v[138] = 10'b1111001111;
    16'b0000100000000011: out_v[138] = 10'b1011011011;
    16'b0100100000000011: out_v[138] = 10'b1100011110;
    16'b0101100000001000: out_v[138] = 10'b0110111110;
    16'b0100000000000010: out_v[138] = 10'b1111111011;
    16'b0100100000000010: out_v[138] = 10'b1111100011;
    16'b0000100000001001: out_v[138] = 10'b0110011000;
    16'b0000110000001000: out_v[138] = 10'b0101010010;
    16'b0000100000011000: out_v[138] = 10'b0110011101;
    16'b0000110000000000: out_v[138] = 10'b0011010010;
    16'b0000010000001000: out_v[138] = 10'b1001010110;
    16'b0000110000100000: out_v[138] = 10'b1111001010;
    16'b0000110000100010: out_v[138] = 10'b1111101100;
    16'b0000110000100011: out_v[138] = 10'b0011001011;
    16'b0000100000011011: out_v[138] = 10'b1110000010;
    16'b0000000000011011: out_v[138] = 10'b1001111110;
    16'b0000100000101001: out_v[138] = 10'b0110011111;
    16'b0000000000101001: out_v[138] = 10'b1011101000;
    16'b0000100000111011: out_v[138] = 10'b1101101011;
    16'b0100100000101010: out_v[138] = 10'b1101010010;
    16'b0000100000101010: out_v[138] = 10'b1101111000;
    16'b0000000000011010: out_v[138] = 10'b1100001111;
    16'b0000100000011010: out_v[138] = 10'b0111110111;
    16'b0000000000010011: out_v[138] = 10'b1010001001;
    default: out_v[138] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100000100100010: out_v[139] = 10'b1100110000;
    16'b1100100100100010: out_v[139] = 10'b0110110011;
    16'b1000100101100110: out_v[139] = 10'b0111001011;
    16'b0100100100100010: out_v[139] = 10'b0010111100;
    16'b1000100101100010: out_v[139] = 10'b1111010001;
    16'b1000100100000110: out_v[139] = 10'b1011010011;
    16'b1000100000100010: out_v[139] = 10'b0101101011;
    16'b1000100100100100: out_v[139] = 10'b0111011101;
    16'b1100100100000010: out_v[139] = 10'b0111100011;
    16'b1100100101100010: out_v[139] = 10'b1000001111;
    16'b1000100100100010: out_v[139] = 10'b1100010011;
    16'b1000100101000010: out_v[139] = 10'b0111000101;
    16'b1000100100100110: out_v[139] = 10'b0010011001;
    16'b0000100100000100: out_v[139] = 10'b1001110011;
    16'b0000100100100010: out_v[139] = 10'b1000110110;
    16'b1000100101100100: out_v[139] = 10'b0110111111;
    16'b0000100100100100: out_v[139] = 10'b1000000011;
    16'b0000100100100110: out_v[139] = 10'b1111001111;
    16'b1000000100100110: out_v[139] = 10'b1001101100;
    16'b1000100100000010: out_v[139] = 10'b0111011011;
    16'b1100100000100010: out_v[139] = 10'b1010111100;
    16'b0000100100000010: out_v[139] = 10'b1100110010;
    16'b1000000100100100: out_v[139] = 10'b1000100100;
    16'b1100100000100000: out_v[139] = 10'b0001011001;
    16'b1100100100100110: out_v[139] = 10'b1000011111;
    16'b0000100100000110: out_v[139] = 10'b1101110111;
    16'b0100000100000010: out_v[139] = 10'b1011100011;
    16'b1100000100100010: out_v[139] = 10'b0111101010;
    16'b1100100101100110: out_v[139] = 10'b1110000011;
    16'b1000000100100010: out_v[139] = 10'b0001111100;
    16'b1000100100000100: out_v[139] = 10'b0110110011;
    16'b0100100100000010: out_v[139] = 10'b0111010100;
    16'b1000000101100110: out_v[139] = 10'b1011000101;
    16'b0100100100100110: out_v[139] = 10'b1001100011;
    16'b1100100101000010: out_v[139] = 10'b1011011000;
    16'b1000000001100000: out_v[139] = 10'b1001011101;
    16'b0000000000100000: out_v[139] = 10'b0001100110;
    16'b0000000100000000: out_v[139] = 10'b0011001101;
    16'b0000000000000000: out_v[139] = 10'b1110000110;
    16'b0000000001000000: out_v[139] = 10'b1010001101;
    16'b0000000100000010: out_v[139] = 10'b0100001110;
    16'b1000000001000000: out_v[139] = 10'b1011011011;
    16'b0000000000000010: out_v[139] = 10'b0110011011;
    16'b1000000000100000: out_v[139] = 10'b1101000111;
    16'b0100000100000000: out_v[139] = 10'b0110111011;
    16'b1100000001000000: out_v[139] = 10'b0011010001;
    16'b1100000000100000: out_v[139] = 10'b1001100011;
    16'b1100000001100000: out_v[139] = 10'b1010010110;
    16'b0000000101000000: out_v[139] = 10'b0010010010;
    16'b1000000000000000: out_v[139] = 10'b0010101111;
    16'b1000000100000000: out_v[139] = 10'b0101001100;
    16'b1100100100100000: out_v[139] = 10'b0010101110;
    16'b1000000101100000: out_v[139] = 10'b0111011101;
    16'b0000000100000100: out_v[139] = 10'b1000100111;
    16'b0100100000000010: out_v[139] = 10'b0111011110;
    16'b1000000100100000: out_v[139] = 10'b0110110100;
    16'b0100100100000000: out_v[139] = 10'b0110100110;
    16'b1100000100000000: out_v[139] = 10'b0010101111;
    16'b0000000000000110: out_v[139] = 10'b0110100100;
    16'b1100100101100000: out_v[139] = 10'b1000111110;
    16'b1000000101100010: out_v[139] = 10'b0011011111;
    16'b0100000100000100: out_v[139] = 10'b0100000010;
    16'b0100100101100000: out_v[139] = 10'b1110100111;
    16'b0000000100100000: out_v[139] = 10'b0110011101;
    16'b1100100100000000: out_v[139] = 10'b1000101110;
    16'b1000100101100000: out_v[139] = 10'b1111011110;
    16'b0000000100000110: out_v[139] = 10'b0011011011;
    16'b1000000100000100: out_v[139] = 10'b0111111010;
    16'b1000000101100100: out_v[139] = 10'b1110101100;
    16'b1100100001100000: out_v[139] = 10'b0010010110;
    16'b1000000100000010: out_v[139] = 10'b1101011110;
    16'b1100100100000100: out_v[139] = 10'b1110010110;
    16'b1100000100100000: out_v[139] = 10'b0000111001;
    16'b1000000100000110: out_v[139] = 10'b0001011100;
    16'b1100000100000100: out_v[139] = 10'b1001011100;
    16'b0000100100000000: out_v[139] = 10'b1111001110;
    16'b1000100100000000: out_v[139] = 10'b0010101010;
    16'b0100000000000110: out_v[139] = 10'b1010001111;
    16'b0000000100100100: out_v[139] = 10'b1010000001;
    16'b1000100001100000: out_v[139] = 10'b0010011110;
    16'b0100100100100000: out_v[139] = 10'b0010101111;
    16'b0100100100000100: out_v[139] = 10'b0011110010;
    16'b1100000101100000: out_v[139] = 10'b1001011010;
    16'b1100000101000000: out_v[139] = 10'b1010100011;
    16'b1100000000000000: out_v[139] = 10'b1100111011;
    16'b0100000100100000: out_v[139] = 10'b0110111110;
    16'b1100000101100010: out_v[139] = 10'b1110000001;
    16'b0100000100100100: out_v[139] = 10'b1101000011;
    16'b1100000100100100: out_v[139] = 10'b1100110011;
    16'b1100000100000110: out_v[139] = 10'b0101011111;
    16'b0100000000000010: out_v[139] = 10'b0011010000;
    16'b0100000000000000: out_v[139] = 10'b0101111100;
    16'b1100000100000010: out_v[139] = 10'b0011111010;
    16'b0100100100000110: out_v[139] = 10'b0110101000;
    16'b0100000100100110: out_v[139] = 10'b0101011011;
    16'b1100000100100110: out_v[139] = 10'b1001101010;
    16'b0100000100000110: out_v[139] = 10'b0101001101;
    16'b0000100000000100: out_v[139] = 10'b0001010010;
    16'b0100100000100000: out_v[139] = 10'b1001010110;
    16'b0000100000100110: out_v[139] = 10'b0110111001;
    16'b0100100000100010: out_v[139] = 10'b1000001101;
    16'b0100100000000100: out_v[139] = 10'b0101010010;
    16'b0000100000100100: out_v[139] = 10'b0001111101;
    16'b0100000000100000: out_v[139] = 10'b0111110010;
    16'b0100100000100100: out_v[139] = 10'b0000011010;
    16'b0100000000000100: out_v[139] = 10'b1100010011;
    16'b0100000000100010: out_v[139] = 10'b1101111101;
    16'b0000100000100010: out_v[139] = 10'b1111000010;
    16'b0100100001000010: out_v[139] = 10'b1000111011;
    16'b0000100000000000: out_v[139] = 10'b1011111001;
    16'b0000100000000010: out_v[139] = 10'b1100011001;
    16'b0000100000100000: out_v[139] = 10'b1011110000;
    16'b0000100001000000: out_v[139] = 10'b1110011001;
    16'b0100100000000000: out_v[139] = 10'b0111010011;
    16'b0100100001100100: out_v[139] = 10'b1010110010;
    16'b0000100001100100: out_v[139] = 10'b1111011010;
    16'b0100100000100110: out_v[139] = 10'b0011111010;
    16'b0100100001000000: out_v[139] = 10'b0110101001;
    16'b0100000000100100: out_v[139] = 10'b1101000111;
    16'b0100100001100010: out_v[139] = 10'b1110011011;
    16'b0100100000000110: out_v[139] = 10'b1110100101;
    16'b1100000000100010: out_v[139] = 10'b1101010000;
    16'b1000000000100010: out_v[139] = 10'b0110010011;
    16'b1000000101000010: out_v[139] = 10'b1110110101;
    16'b1000000101000100: out_v[139] = 10'b0011100010;
    16'b1100000101000010: out_v[139] = 10'b0010110000;
    16'b1100000000000010: out_v[139] = 10'b1100100010;
    16'b0100000101000010: out_v[139] = 10'b1001111000;
    16'b1100000000100110: out_v[139] = 10'b0100011011;
    16'b0100100100100100: out_v[139] = 10'b1111000111;
    16'b0000100101000010: out_v[139] = 10'b0001110001;
    16'b0100100101000010: out_v[139] = 10'b0011010110;
    16'b0100000101000000: out_v[139] = 10'b0111000110;
    16'b0100000001000000: out_v[139] = 10'b0101010000;
    16'b0000100000000110: out_v[139] = 10'b0110000011;
    16'b1100100001000000: out_v[139] = 10'b1011000111;
    16'b0100100101000000: out_v[139] = 10'b1011000000;
    16'b0000000000000100: out_v[139] = 10'b1101110000;
    16'b0000000000100110: out_v[139] = 10'b0010100000;
    16'b0000000000100010: out_v[139] = 10'b0011001100;
    16'b0000000000100100: out_v[139] = 10'b0110000101;
    16'b0000010000000110: out_v[139] = 10'b0011111011;
    16'b0000000100100110: out_v[139] = 10'b0111001010;
    16'b0000010000100110: out_v[139] = 10'b1110110101;
    16'b0000000100100010: out_v[139] = 10'b0111111001;
    16'b0000000000010110: out_v[139] = 10'b1110110010;
    16'b0000000000110110: out_v[139] = 10'b0100110111;
    16'b1000000000100110: out_v[139] = 10'b1000010110;
    16'b1100100100100100: out_v[139] = 10'b0110000110;
    16'b0100000101100010: out_v[139] = 10'b1111001010;
    16'b0100000000100110: out_v[139] = 10'b1100101110;
    default: out_v[139] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1001000110100000: out_v[140] = 10'b1101110001;
    16'b1101000110100000: out_v[140] = 10'b0010001111;
    16'b1101000100100100: out_v[140] = 10'b1111101110;
    16'b0101000100100100: out_v[140] = 10'b0111111011;
    16'b1101000110000000: out_v[140] = 10'b0100011010;
    16'b1101000000000100: out_v[140] = 10'b1000011011;
    16'b1101000110000100: out_v[140] = 10'b1001001011;
    16'b0101000000100100: out_v[140] = 10'b1101010011;
    16'b0100000000000100: out_v[140] = 10'b1101011011;
    16'b0110100100100000: out_v[140] = 10'b0111001011;
    16'b1101001110100000: out_v[140] = 10'b0011100101;
    16'b0111100100100000: out_v[140] = 10'b1011001011;
    16'b0101000110100000: out_v[140] = 10'b0100100011;
    16'b1101000010000100: out_v[140] = 10'b1101010011;
    16'b1001000110000000: out_v[140] = 10'b1111000111;
    16'b1001100110100000: out_v[140] = 10'b1010110011;
    16'b1111000110100100: out_v[140] = 10'b1110110000;
    16'b0101100100100000: out_v[140] = 10'b1010010001;
    16'b1101000110100100: out_v[140] = 10'b0000001111;
    16'b1001000110100100: out_v[140] = 10'b0111111001;
    16'b0100000100100100: out_v[140] = 10'b0110110010;
    16'b0100000000100100: out_v[140] = 10'b0101110001;
    16'b0101100100100100: out_v[140] = 10'b0111110011;
    16'b0110000000100100: out_v[140] = 10'b0101010011;
    16'b0100100100100000: out_v[140] = 10'b1011011111;
    16'b1000000110100000: out_v[140] = 10'b1001011001;
    16'b0110000100100000: out_v[140] = 10'b1100110110;
    16'b0101000100000100: out_v[140] = 10'b1010010000;
    16'b0101000100100000: out_v[140] = 10'b1101110011;
    16'b1101001110100100: out_v[140] = 10'b1110010101;
    16'b0110100100000000: out_v[140] = 10'b0011011011;
    16'b1000000010100000: out_v[140] = 10'b0110100101;
    16'b0101100100000000: out_v[140] = 10'b1001110001;
    16'b1001000110000100: out_v[140] = 10'b1111100011;
    16'b1111000110100000: out_v[140] = 10'b1000011101;
    16'b0100000100100000: out_v[140] = 10'b1100110001;
    16'b0101000100000000: out_v[140] = 10'b1001001010;
    16'b1000000110000000: out_v[140] = 10'b0011010000;
    16'b1101100110100000: out_v[140] = 10'b0011111010;
    16'b0101000000000100: out_v[140] = 10'b1101101011;
    16'b0111000100100100: out_v[140] = 10'b0101010101;
    16'b0110000100100100: out_v[140] = 10'b1111111110;
    16'b1001000010100000: out_v[140] = 10'b0110100110;
    16'b0111000100100000: out_v[140] = 10'b1101011111;
    16'b0110000100000000: out_v[140] = 10'b0110111001;
    16'b1101001110000100: out_v[140] = 10'b0111010111;
    16'b0110100000100100: out_v[140] = 10'b1011011110;
    16'b0000001000100000: out_v[140] = 10'b0010001010;
    16'b0000001000000000: out_v[140] = 10'b0011100011;
    16'b0000000000000000: out_v[140] = 10'b0011001100;
    16'b1000000000000000: out_v[140] = 10'b1001011001;
    16'b0000000000100000: out_v[140] = 10'b0010100111;
    16'b1000100000000000: out_v[140] = 10'b1110011011;
    16'b1000001000000000: out_v[140] = 10'b1100011101;
    16'b1000001000100000: out_v[140] = 10'b1100010010;
    16'b0000100000000000: out_v[140] = 10'b0000010110;
    16'b1000101000000000: out_v[140] = 10'b0001110010;
    16'b1000000010000000: out_v[140] = 10'b1101010010;
    16'b1000000000100000: out_v[140] = 10'b0110100001;
    16'b0010101000000000: out_v[140] = 10'b1111001101;
    16'b0000100100000100: out_v[140] = 10'b1011100100;
    16'b0000101000100000: out_v[140] = 10'b1101111101;
    16'b0010101000100000: out_v[140] = 10'b0011000101;
    16'b0000100100000000: out_v[140] = 10'b1000001000;
    16'b0000000100000000: out_v[140] = 10'b0010111100;
    16'b0010001000000000: out_v[140] = 10'b0001011110;
    16'b0000100000100000: out_v[140] = 10'b0001011010;
    16'b0010100100000000: out_v[140] = 10'b1011011011;
    16'b0000001100000100: out_v[140] = 10'b0101100100;
    16'b0010101100000000: out_v[140] = 10'b0011101000;
    16'b0010000000000000: out_v[140] = 10'b1101110111;
    16'b0010100100000100: out_v[140] = 10'b1000001011;
    16'b0010000100000100: out_v[140] = 10'b0001100001;
    16'b0000101000000000: out_v[140] = 10'b1101100101;
    16'b0000000100000100: out_v[140] = 10'b0000100110;
    16'b0000100100100100: out_v[140] = 10'b1010010110;
    16'b0000101100000000: out_v[140] = 10'b1010101110;
    16'b0000001100000000: out_v[140] = 10'b0110100010;
    16'b0000100000000100: out_v[140] = 10'b1001010101;
    16'b0010100000000000: out_v[140] = 10'b0010110101;
    16'b0010100000100000: out_v[140] = 10'b1110111010;
    16'b0000101100000100: out_v[140] = 10'b1010110011;
    16'b0010101100000100: out_v[140] = 10'b1011100101;
    16'b0000000000000100: out_v[140] = 10'b0111001000;
    16'b0000100100100000: out_v[140] = 10'b1011010110;
    16'b0010001000100000: out_v[140] = 10'b1001111110;
    16'b0010000000100000: out_v[140] = 10'b0000001110;
    16'b1000001010100000: out_v[140] = 10'b0110010111;
    16'b0000101010100000: out_v[140] = 10'b1101110101;
    16'b1010000010100000: out_v[140] = 10'b1011111001;
    16'b1000101010100000: out_v[140] = 10'b0011011000;
    16'b0000001100100000: out_v[140] = 10'b0010001001;
    16'b0000001010100000: out_v[140] = 10'b0010001101;
    16'b1111000010100000: out_v[140] = 10'b0001110110;
    16'b1000001010000000: out_v[140] = 10'b1110110000;
    16'b1000101000100000: out_v[140] = 10'b1111000011;
    16'b0000001000100100: out_v[140] = 10'b1111111001;
    16'b0010001100100000: out_v[140] = 10'b1011110011;
    16'b1001101010100000: out_v[140] = 10'b1111010111;
    16'b1111001010100000: out_v[140] = 10'b1110111010;
    16'b1010001010100000: out_v[140] = 10'b1010011111;
    16'b0000001000000100: out_v[140] = 10'b1000001001;
    16'b1000101010100100: out_v[140] = 10'b0011010111;
    16'b0000101000100100: out_v[140] = 10'b1011110011;
    16'b1000001110100000: out_v[140] = 10'b1001001010;
    16'b1111101010100000: out_v[140] = 10'b1001111011;
    16'b0010001010100000: out_v[140] = 10'b1011110111;
    16'b1000001010100100: out_v[140] = 10'b1011011111;
    16'b1100001010100000: out_v[140] = 10'b0000111110;
    16'b1001001010100000: out_v[140] = 10'b1101010100;
    16'b1101101010100000: out_v[140] = 10'b0001001010;
    16'b1101100010100000: out_v[140] = 10'b1010111101;
    16'b1000101010000000: out_v[140] = 10'b0011101011;
    16'b0000000000100100: out_v[140] = 10'b0011111001;
    16'b1000100010100000: out_v[140] = 10'b1001001111;
    16'b0000000100100000: out_v[140] = 10'b0010001110;
    16'b1101001010100000: out_v[140] = 10'b0011101110;
    16'b1000100000100000: out_v[140] = 10'b1110011001;
    16'b0100001100000000: out_v[140] = 10'b1000010000;
    16'b0101000010100000: out_v[140] = 10'b1100110101;
    16'b0101001100000000: out_v[140] = 10'b0101010010;
    16'b0101001100100000: out_v[140] = 10'b1000010111;
    16'b0100000000000000: out_v[140] = 10'b1000111010;
    16'b0100000100000000: out_v[140] = 10'b1100011011;
    16'b0100001000000000: out_v[140] = 10'b1101011111;
    16'b1001001110100000: out_v[140] = 10'b0101100111;
    16'b1101000010100000: out_v[140] = 10'b0010111010;
    16'b0101000000000000: out_v[140] = 10'b1100111100;
    16'b1001001010000000: out_v[140] = 10'b1001110110;
    16'b1101001110000000: out_v[140] = 10'b0011101110;
    16'b0111000100000000: out_v[140] = 10'b0001010011;
    16'b0110001100000000: out_v[140] = 10'b1110011011;
    16'b1001001110000000: out_v[140] = 10'b0101011011;
    16'b0101000010000000: out_v[140] = 10'b0110100110;
    16'b0101000000100000: out_v[140] = 10'b1111000010;
    16'b0101001000000000: out_v[140] = 10'b0011010110;
    16'b0101000110000000: out_v[140] = 10'b0010101001;
    16'b1101000100000000: out_v[140] = 10'b1100001001;
    16'b0010000100000000: out_v[140] = 10'b1110000111;
    16'b1101000010000000: out_v[140] = 10'b0010010100;
    16'b1000001110000000: out_v[140] = 10'b0101110001;
    16'b0001001000000000: out_v[140] = 10'b1001100001;
    16'b0100000100000100: out_v[140] = 10'b1001111011;
    16'b0101001010000000: out_v[140] = 10'b0101111001;
    16'b1001000010000000: out_v[140] = 10'b1010000111;
    16'b0101001110000000: out_v[140] = 10'b0011101101;
    16'b0001001010000000: out_v[140] = 10'b0101011001;
    16'b1101001010000000: out_v[140] = 10'b0110100110;
    16'b0001000010100000: out_v[140] = 10'b1101010010;
    16'b1000001010000100: out_v[140] = 10'b1010001100;
    16'b0100000000100000: out_v[140] = 10'b1101100010;
    16'b1001000010100100: out_v[140] = 10'b1111011111;
    16'b1001000010000100: out_v[140] = 10'b1110110001;
    16'b1101000010100100: out_v[140] = 10'b1000011100;
    16'b0111000010100000: out_v[140] = 10'b0111110001;
    16'b1000000010000100: out_v[140] = 10'b1110000010;
    16'b0001000010000000: out_v[140] = 10'b1101110001;
    16'b1001100010100000: out_v[140] = 10'b0101110011;
    16'b0100000010100000: out_v[140] = 10'b1101100010;
    16'b0110000010100000: out_v[140] = 10'b0111100010;
    16'b0110000000100000: out_v[140] = 10'b0111010111;
    16'b1111000110000000: out_v[140] = 10'b1110011101;
    16'b0101100100010000: out_v[140] = 10'b1011101111;
    16'b0101100110000000: out_v[140] = 10'b1111101011;
    16'b0100100100000000: out_v[140] = 10'b0111010011;
    16'b1000100010010000: out_v[140] = 10'b1111000010;
    16'b1101100110010000: out_v[140] = 10'b0111101000;
    16'b1001100010000000: out_v[140] = 10'b1110111000;
    16'b1001100010010000: out_v[140] = 10'b1010100011;
    16'b0100101100000000: out_v[140] = 10'b1011011000;
    16'b1101100110000000: out_v[140] = 10'b1011011100;
    16'b1101101110000000: out_v[140] = 10'b1011000110;
    16'b1001100110010000: out_v[140] = 10'b1110110100;
    16'b0100100100010000: out_v[140] = 10'b0111111011;
    16'b0111100100000000: out_v[140] = 10'b0001011100;
    16'b0101100110010000: out_v[140] = 10'b1100011111;
    16'b0001100010010000: out_v[140] = 10'b0001011011;
    16'b0101101100000000: out_v[140] = 10'b1011011011;
    16'b1101000000100000: out_v[140] = 10'b0101010011;
    16'b1001000000100000: out_v[140] = 10'b0011011100;
    16'b1001001000000000: out_v[140] = 10'b0011100010;
    16'b1101000000000000: out_v[140] = 10'b1010000100;
    16'b0001000000100000: out_v[140] = 10'b0101111110;
    16'b1101001000000000: out_v[140] = 10'b0101100100;
    16'b1001000000000000: out_v[140] = 10'b1111001010;
    16'b1001001000100000: out_v[140] = 10'b1011011001;
    16'b1101001000100000: out_v[140] = 10'b1101001010;
    16'b0001000000000000: out_v[140] = 10'b1111100000;
    16'b0101001000100000: out_v[140] = 10'b0010011110;
    16'b1000000100100000: out_v[140] = 10'b0111101100;
    16'b1000001100100000: out_v[140] = 10'b1100010110;
    16'b0001001010100000: out_v[140] = 10'b1101010001;
    16'b0101001010100000: out_v[140] = 10'b1100000010;
    16'b0100001101000000: out_v[140] = 10'b1001110101;
    16'b0100000101000000: out_v[140] = 10'b0111011010;
    16'b0101001101000000: out_v[140] = 10'b0111001111;
    16'b1101000100100000: out_v[140] = 10'b1100001001;
    16'b0110000101000000: out_v[140] = 10'b0001100101;
    16'b0100001001000000: out_v[140] = 10'b1110000101;
    16'b0101001001000000: out_v[140] = 10'b1111100001;
    16'b1101001100000000: out_v[140] = 10'b1000100011;
    16'b0000000101000000: out_v[140] = 10'b1001100111;
    16'b0101000101000000: out_v[140] = 10'b0111100111;
    default: out_v[140] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010001000111010: out_v[141] = 10'b0000111011;
    16'b0001001000001000: out_v[141] = 10'b0110010011;
    16'b0011001000111010: out_v[141] = 10'b1100011110;
    16'b0010001000011010: out_v[141] = 10'b1000100110;
    16'b0111001000111010: out_v[141] = 10'b1011110110;
    16'b0000001000011000: out_v[141] = 10'b1110010001;
    16'b0000001000001000: out_v[141] = 10'b0010100111;
    16'b0001001000011000: out_v[141] = 10'b1111101010;
    16'b0001001000011010: out_v[141] = 10'b1011111100;
    16'b0001000000011000: out_v[141] = 10'b1110111101;
    16'b0010001000110010: out_v[141] = 10'b1000010001;
    16'b0110001000111010: out_v[141] = 10'b1010010011;
    16'b0011000000011000: out_v[141] = 10'b1011111011;
    16'b0001001000101010: out_v[141] = 10'b0000000011;
    16'b0011001000011000: out_v[141] = 10'b0111111001;
    16'b0010001000011000: out_v[141] = 10'b0110010111;
    16'b0011001000011010: out_v[141] = 10'b1101111110;
    16'b0001001000100010: out_v[141] = 10'b1010111111;
    16'b0011001000110010: out_v[141] = 10'b0011001101;
    16'b0001001000111010: out_v[141] = 10'b0011000111;
    16'b0011000000011010: out_v[141] = 10'b0100001110;
    16'b0000011000011000: out_v[141] = 10'b1111000010;
    16'b0011000000111010: out_v[141] = 10'b1110010011;
    16'b0000001000010000: out_v[141] = 10'b0110001111;
    16'b0010000000111010: out_v[141] = 10'b0000100000;
    16'b0000001000000000: out_v[141] = 10'b0000010101;
    16'b0110011000111010: out_v[141] = 10'b0010001011;
    16'b0000001000011010: out_v[141] = 10'b1110010011;
    16'b0110010000111010: out_v[141] = 10'b1011110111;
    16'b0000001000111010: out_v[141] = 10'b1110010001;
    16'b0100010001000100: out_v[141] = 10'b0010010010;
    16'b0000000001000100: out_v[141] = 10'b1100110110;
    16'b0100000001000000: out_v[141] = 10'b1110111001;
    16'b0000000001000000: out_v[141] = 10'b1001000011;
    16'b0000000000000000: out_v[141] = 10'b0000111001;
    16'b0100010001000000: out_v[141] = 10'b0100100001;
    16'b0100000001000100: out_v[141] = 10'b1101101000;
    16'b0100011001000100: out_v[141] = 10'b0110011000;
    16'b0100011001000000: out_v[141] = 10'b1100011010;
    16'b0100011001000101: out_v[141] = 10'b1000011010;
    16'b0010000001000100: out_v[141] = 10'b0011000001;
    16'b0000010001000100: out_v[141] = 10'b0001001001;
    16'b0000000001000110: out_v[141] = 10'b1010010011;
    16'b0100010001100110: out_v[141] = 10'b1101010101;
    16'b0100010001101110: out_v[141] = 10'b0100110001;
    16'b0100010001001110: out_v[141] = 10'b0111110100;
    16'b0100010001101010: out_v[141] = 10'b1110001101;
    16'b0100010001001000: out_v[141] = 10'b1110000110;
    16'b0000011001001100: out_v[141] = 10'b0110110111;
    16'b0110010001010100: out_v[141] = 10'b0000110100;
    16'b0110010001111110: out_v[141] = 10'b1001001111;
    16'b0110011001101110: out_v[141] = 10'b0010110111;
    16'b0110011001001100: out_v[141] = 10'b1001100111;
    16'b0000001001001000: out_v[141] = 10'b0110000111;
    16'b0100011001101110: out_v[141] = 10'b1100000111;
    16'b0100010001000110: out_v[141] = 10'b1101010100;
    16'b0000011001000100: out_v[141] = 10'b1100001101;
    16'b0100011001001100: out_v[141] = 10'b1111101100;
    16'b0110010001011100: out_v[141] = 10'b0011000100;
    16'b0100010001001100: out_v[141] = 10'b1000110100;
    16'b0110010001001100: out_v[141] = 10'b0111100101;
    16'b0010011001001100: out_v[141] = 10'b1110101011;
    16'b0000011001101110: out_v[141] = 10'b0110110010;
    16'b0110011001011100: out_v[141] = 10'b1000011100;
    16'b0000011001100110: out_v[141] = 10'b0100100110;
    16'b0110011001111110: out_v[141] = 10'b0110010101;
    16'b0100000001101110: out_v[141] = 10'b1010111101;
    16'b0000000001101110: out_v[141] = 10'b1101001001;
    16'b0110010001011110: out_v[141] = 10'b1100100101;
    16'b0000000001100110: out_v[141] = 10'b1111010100;
    16'b0100010000000000: out_v[141] = 10'b1010110111;
    16'b0110010001000100: out_v[141] = 10'b1011101011;
    16'b0010011001011100: out_v[141] = 10'b0000110111;
    16'b0100011001100110: out_v[141] = 10'b1001101101;
    16'b0100011001001110: out_v[141] = 10'b1110011011;
    16'b0110010001101110: out_v[141] = 10'b1110100110;
    16'b0010011001111110: out_v[141] = 10'b0000101100;
    16'b0000011001001110: out_v[141] = 10'b1100111111;
    16'b0000000001001100: out_v[141] = 10'b1111000101;
    16'b0100011001101010: out_v[141] = 10'b1111101111;
    16'b0000001001001100: out_v[141] = 10'b1000110110;
    16'b0010000001001100: out_v[141] = 10'b1010010110;
    16'b0100010000101010: out_v[141] = 10'b1010011011;
    16'b0000000000001010: out_v[141] = 10'b1111000010;
    16'b0100010000001000: out_v[141] = 10'b0111100111;
    16'b0100011000001010: out_v[141] = 10'b1111001011;
    16'b0100010000111010: out_v[141] = 10'b1111011010;
    16'b0000010000101010: out_v[141] = 10'b1011101010;
    16'b0010010000101010: out_v[141] = 10'b1101001011;
    16'b0100011000101010: out_v[141] = 10'b1001001001;
    16'b0110010000001000: out_v[141] = 10'b1101011110;
    16'b0100010000100010: out_v[141] = 10'b1011001110;
    16'b0110011000001000: out_v[141] = 10'b0101011010;
    16'b0000000000001000: out_v[141] = 10'b1011000111;
    16'b0100011000001000: out_v[141] = 10'b1100000011;
    16'b0000010000100010: out_v[141] = 10'b1101010100;
    16'b0100000000001010: out_v[141] = 10'b1111010101;
    16'b0100010000001010: out_v[141] = 10'b0010111011;
    16'b0100000000101010: out_v[141] = 10'b0001011110;
    16'b0110011000011000: out_v[141] = 10'b0001011100;
    16'b0100011000101011: out_v[141] = 10'b1101111111;
    16'b0000000000101010: out_v[141] = 10'b1011001110;
    16'b0110010000101010: out_v[141] = 10'b1001001100;
    16'b0000010000001010: out_v[141] = 10'b0011111101;
    16'b0110011000001010: out_v[141] = 10'b1001111011;
    16'b0000000000100010: out_v[141] = 10'b0010110111;
    16'b0100011000000000: out_v[141] = 10'b0100011010;
    16'b0000010000000000: out_v[141] = 10'b0011101100;
    16'b0000010000001000: out_v[141] = 10'b1111100100;
    16'b0110011000101010: out_v[141] = 10'b0111001011;
    16'b0000010000110010: out_v[141] = 10'b0100110110;
    16'b0110010000001010: out_v[141] = 10'b1010111101;
    16'b0100000000001000: out_v[141] = 10'b0001010110;
    16'b0100000000000000: out_v[141] = 10'b1110101000;
    16'b0000010000111010: out_v[141] = 10'b0011011101;
    16'b0110010000100010: out_v[141] = 10'b0000011000;
    16'b0010010000111010: out_v[141] = 10'b1010100110;
    16'b0100010001111110: out_v[141] = 10'b0100110011;
    16'b0010011000010000: out_v[141] = 10'b0001111111;
    16'b0010011001010100: out_v[141] = 10'b0101110011;
    16'b0110011001010100: out_v[141] = 10'b0011011010;
    16'b0110011001010000: out_v[141] = 10'b1000011111;
    16'b0100010001010100: out_v[141] = 10'b0000011011;
    16'b0000011001010100: out_v[141] = 10'b0100011011;
    16'b0100011001010000: out_v[141] = 10'b0111000111;
    16'b0110010001010000: out_v[141] = 10'b1001011110;
    16'b0100011000010000: out_v[141] = 10'b1111000010;
    16'b0110010001111010: out_v[141] = 10'b1010101110;
    16'b0100010001010000: out_v[141] = 10'b1101100110;
    16'b0100011001010100: out_v[141] = 10'b1011000111;
    16'b0100010000010000: out_v[141] = 10'b1110000101;
    16'b0110011000010000: out_v[141] = 10'b1010011010;
    16'b0100010001111010: out_v[141] = 10'b0111010000;
    16'b0110010000010000: out_v[141] = 10'b1011000110;
    16'b0100010001001010: out_v[141] = 10'b1111110100;
    16'b0000011000000000: out_v[141] = 10'b1110010111;
    16'b0010011001010000: out_v[141] = 10'b1001000111;
    16'b0000011000010000: out_v[141] = 10'b0011011011;
    16'b0000011001010000: out_v[141] = 10'b0100011010;
    16'b0100010001011010: out_v[141] = 10'b0100110111;
    16'b0100001000000000: out_v[141] = 10'b1111100010;
    16'b0010010000011010: out_v[141] = 10'b1001100010;
    16'b0100001001000100: out_v[141] = 10'b0001101100;
    16'b0000000001010100: out_v[141] = 10'b0010011110;
    16'b0000000000111010: out_v[141] = 10'b1101110110;
    16'b0000000000010000: out_v[141] = 10'b0110111111;
    16'b0000010000011000: out_v[141] = 10'b0101111101;
    16'b0100001001010100: out_v[141] = 10'b1111100101;
    16'b0000000000011000: out_v[141] = 10'b1111001011;
    16'b0010010000110010: out_v[141] = 10'b0001110010;
    16'b0010000000010000: out_v[141] = 10'b1101100101;
    16'b0010000000011000: out_v[141] = 10'b0101010111;
    16'b0010000001010100: out_v[141] = 10'b1100110101;
    16'b0000010000011010: out_v[141] = 10'b1011011100;
    16'b0010000000011010: out_v[141] = 10'b0001011001;
    16'b0000010000010000: out_v[141] = 10'b0100111000;
    16'b0000001001010100: out_v[141] = 10'b1101001111;
    16'b0000001001000100: out_v[141] = 10'b0101110100;
    16'b0000000001010000: out_v[141] = 10'b0000101100;
    16'b0100010000110010: out_v[141] = 10'b0100010110;
    16'b0010010000011000: out_v[141] = 10'b0101110110;
    16'b0010000001111110: out_v[141] = 10'b0101001010;
    16'b0010000001111010: out_v[141] = 10'b1010011011;
    16'b0110010000110010: out_v[141] = 10'b0110100010;
    16'b0010000001010000: out_v[141] = 10'b0010111111;
    16'b0000000000011010: out_v[141] = 10'b1101001101;
    16'b0010000001011010: out_v[141] = 10'b1000111110;
    16'b0110010000011010: out_v[141] = 10'b1001110101;
    16'b0000000001011100: out_v[141] = 10'b1101000111;
    16'b0010010001111110: out_v[141] = 10'b0101011010;
    16'b0000010001011000: out_v[141] = 10'b1010111011;
    16'b0010010001011000: out_v[141] = 10'b1101010010;
    16'b0000010001111110: out_v[141] = 10'b1011000111;
    16'b0010010001011100: out_v[141] = 10'b1101101011;
    16'b0000010001001100: out_v[141] = 10'b1011100101;
    16'b0000010001011100: out_v[141] = 10'b1001101011;
    16'b0000010001001110: out_v[141] = 10'b1000111101;
    16'b0010010001011110: out_v[141] = 10'b1100100111;
    16'b0000000001001110: out_v[141] = 10'b1001110101;
    16'b0000000001011110: out_v[141] = 10'b1111000011;
    16'b0000010001011110: out_v[141] = 10'b1110001001;
    16'b0000000001111110: out_v[141] = 10'b0111000011;
    16'b0000000001001000: out_v[141] = 10'b1111001011;
    16'b0000000001001010: out_v[141] = 10'b1011101001;
    16'b0011010001011100: out_v[141] = 10'b0110111101;
    16'b0100010001011100: out_v[141] = 10'b1000111001;
    16'b0000010001011010: out_v[141] = 10'b1111000110;
    16'b0000010001001000: out_v[141] = 10'b1001100111;
    16'b0010010001111010: out_v[141] = 10'b0001101010;
    16'b0010010001011010: out_v[141] = 10'b1110011110;
    16'b0010000001011110: out_v[141] = 10'b0111100010;
    16'b0111011001011110: out_v[141] = 10'b1011101011;
    16'b0111011001011100: out_v[141] = 10'b0010011101;
    16'b0000010001000000: out_v[141] = 10'b1100011100;
    16'b0010000001011100: out_v[141] = 10'b0010101101;
    16'b0100011000011000: out_v[141] = 10'b0111001111;
    16'b0110010000011000: out_v[141] = 10'b1100110001;
    16'b0100011000010100: out_v[141] = 10'b0101010010;
    16'b0110010000000000: out_v[141] = 10'b0111111111;
    16'b0100001000111010: out_v[141] = 10'b0000100111;
    16'b0010001000010000: out_v[141] = 10'b0011111001;
    16'b0110011000010100: out_v[141] = 10'b0011111101;
    16'b0110011001010101: out_v[141] = 10'b0110110011;
    16'b0110011001000100: out_v[141] = 10'b0111110001;
    16'b0110011000011010: out_v[141] = 10'b0101011100;
    16'b0010011000010100: out_v[141] = 10'b1001011111;
    16'b0010011001000100: out_v[141] = 10'b0111110110;
    16'b0010011000011000: out_v[141] = 10'b1001000111;
    16'b0010011000000000: out_v[141] = 10'b1100100111;
    16'b0010011001010101: out_v[141] = 10'b0100110110;
    16'b0100011000111010: out_v[141] = 10'b0110001101;
    16'b0110011000000000: out_v[141] = 10'b0001101011;
    16'b0000011001010101: out_v[141] = 10'b0011101100;
    16'b0110010001000000: out_v[141] = 10'b1111110010;
    16'b0110011001011110: out_v[141] = 10'b1110011000;
    16'b0110011001111010: out_v[141] = 10'b1110011000;
    16'b0010011001111010: out_v[141] = 10'b1110010000;
    16'b0100011001111010: out_v[141] = 10'b1011101011;
    16'b0110011001011000: out_v[141] = 10'b0110111011;
    16'b0100011001111110: out_v[141] = 10'b1010011001;
    16'b0110011001011010: out_v[141] = 10'b1010011011;
    16'b0011011001010100: out_v[141] = 10'b1010100110;
    16'b0110010001011010: out_v[141] = 10'b1011000111;
    16'b0010010000010000: out_v[141] = 10'b0000110101;
    default: out_v[141] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001000010000100: out_v[142] = 10'b1110100100;
    16'b0001000010000111: out_v[142] = 10'b1011101111;
    16'b0001000000000101: out_v[142] = 10'b1101010001;
    16'b0001000000000001: out_v[142] = 10'b0000100011;
    16'b0101000001000100: out_v[142] = 10'b1010001100;
    16'b0001000011000101: out_v[142] = 10'b1000110011;
    16'b0000000000000101: out_v[142] = 10'b0110010011;
    16'b0001000000000100: out_v[142] = 10'b0111011001;
    16'b0000000000000001: out_v[142] = 10'b1101000001;
    16'b0001000010000101: out_v[142] = 10'b0001001011;
    16'b0101000011000100: out_v[142] = 10'b1100100011;
    16'b0001000001000101: out_v[142] = 10'b0111100010;
    16'b0000000001000101: out_v[142] = 10'b1010100110;
    16'b0101000000000101: out_v[142] = 10'b1111001111;
    16'b0001000000000000: out_v[142] = 10'b0010100111;
    16'b0001000000000111: out_v[142] = 10'b0111010011;
    16'b0101000011000101: out_v[142] = 10'b0101011010;
    16'b0001000010000001: out_v[142] = 10'b1011100010;
    16'b0000000000000100: out_v[142] = 10'b1011110001;
    16'b0001000011000001: out_v[142] = 10'b0101010110;
    16'b0101000000000100: out_v[142] = 10'b0001111101;
    16'b0101000001000101: out_v[142] = 10'b0101000110;
    16'b0101000010000100: out_v[142] = 10'b0111110000;
    16'b0000000000000000: out_v[142] = 10'b1000100111;
    16'b0001000001000001: out_v[142] = 10'b0110000111;
    16'b0101000010000101: out_v[142] = 10'b0100000010;
    16'b0101000010000000: out_v[142] = 10'b0100101000;
    16'b0101000000000000: out_v[142] = 10'b1001101101;
    16'b0000000010000000: out_v[142] = 10'b1100000110;
    16'b0000000010000100: out_v[142] = 10'b1010001110;
    16'b0000000001000100: out_v[142] = 10'b1101100110;
    16'b0000000011000100: out_v[142] = 10'b0101101100;
    16'b0100000011000100: out_v[142] = 10'b0000010111;
    16'b0001000010000000: out_v[142] = 10'b0100011110;
    16'b0100000000000000: out_v[142] = 10'b1010110000;
    16'b0100000010000000: out_v[142] = 10'b0001110000;
    16'b0101000000000010: out_v[142] = 10'b0101100111;
    16'b0000000001000000: out_v[142] = 10'b1011110000;
    16'b0101000011000000: out_v[142] = 10'b0101001111;
    16'b0100000001000000: out_v[142] = 10'b1000010110;
    16'b0000000001000001: out_v[142] = 10'b0000011110;
    16'b0101000001000000: out_v[142] = 10'b1011000110;
    16'b0100000000000100: out_v[142] = 10'b1001001101;
    16'b0001000001000000: out_v[142] = 10'b0110111111;
    16'b0101000011000001: out_v[142] = 10'b0110110101;
    16'b0100000011000001: out_v[142] = 10'b0010011110;
    16'b0100000001000100: out_v[142] = 10'b0010000111;
    16'b0100000011000000: out_v[142] = 10'b0001110111;
    16'b0100000001000001: out_v[142] = 10'b1001001010;
    16'b0000000011000000: out_v[142] = 10'b0111001101;
    16'b0101000001000001: out_v[142] = 10'b1011001000;
    16'b0100000010000100: out_v[142] = 10'b1000101101;
    16'b0100000001000101: out_v[142] = 10'b1010010010;
    16'b0101000000000001: out_v[142] = 10'b1001001111;
    16'b0100000000000101: out_v[142] = 10'b0111010000;
    16'b0001000011000000: out_v[142] = 10'b0001001000;
    16'b0100000011000101: out_v[142] = 10'b1001011100;
    16'b0100000000000001: out_v[142] = 10'b1011010110;
    16'b0101000010000001: out_v[142] = 10'b0110001000;
    16'b0100000010000010: out_v[142] = 10'b0011011010;
    16'b0101000010000010: out_v[142] = 10'b1000000101;
    16'b0001000011000100: out_v[142] = 10'b0111010010;
    16'b0101000010000111: out_v[142] = 10'b0001111011;
    16'b0101000011000110: out_v[142] = 10'b1000110110;
    16'b0001000011000010: out_v[142] = 10'b1110011011;
    16'b0101000010000110: out_v[142] = 10'b0100010100;
    16'b0101001010000100: out_v[142] = 10'b0001111111;
    16'b0101000011000010: out_v[142] = 10'b0100010111;
    16'b0101000011000111: out_v[142] = 10'b1111000110;
    16'b0001000010000010: out_v[142] = 10'b1011100101;
    16'b0100000010000001: out_v[142] = 10'b1100010010;
    16'b0001000011100101: out_v[142] = 10'b1011111110;
    16'b0001000011100100: out_v[142] = 10'b1101011110;
    16'b0000000011100001: out_v[142] = 10'b0111011111;
    16'b0001000001100100: out_v[142] = 10'b1101100111;
    16'b0001000001000100: out_v[142] = 10'b0111010011;
    16'b0001000011000110: out_v[142] = 10'b1110010111;
    16'b0001000011100000: out_v[142] = 10'b0010011011;
    16'b0001000010100100: out_v[142] = 10'b1000110101;
    16'b0000000010000001: out_v[142] = 10'b0001110000;
    16'b0000000011000001: out_v[142] = 10'b1010110110;
    16'b0001000010100001: out_v[142] = 10'b1010111111;
    16'b1001000010000000: out_v[142] = 10'b1111011010;
    16'b1001000011000000: out_v[142] = 10'b1101100010;
    16'b1101000011000000: out_v[142] = 10'b1011010000;
    16'b1101000010000100: out_v[142] = 10'b1011011111;
    16'b1100000011000100: out_v[142] = 10'b1110010101;
    16'b1100000011000000: out_v[142] = 10'b0111100110;
    16'b0100001001000100: out_v[142] = 10'b0011111000;
    16'b0100001001000000: out_v[142] = 10'b1011100010;
    16'b0100001000000100: out_v[142] = 10'b1111100111;
    16'b0100001001000001: out_v[142] = 10'b1001101011;
    16'b0101000000000111: out_v[142] = 10'b0010011111;
    16'b0101000000000110: out_v[142] = 10'b0011111011;
    16'b0101000001000111: out_v[142] = 10'b0011100011;
    16'b0000001001000101: out_v[142] = 10'b1100100011;
    16'b0100001001000101: out_v[142] = 10'b1111010000;
    16'b0101001001000101: out_v[142] = 10'b1101100111;
    16'b0101000001000110: out_v[142] = 10'b0011111010;
    16'b0101000011100101: out_v[142] = 10'b1011001110;
    16'b0101000010100101: out_v[142] = 10'b1001011111;
    16'b0100000010000101: out_v[142] = 10'b0110001110;
    16'b0100000010000111: out_v[142] = 10'b1001001110;
    default: out_v[142] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000010100001001: out_v[143] = 10'b1000110111;
    16'b1100010000000101: out_v[143] = 10'b0000000111;
    16'b1100010100000001: out_v[143] = 10'b0100100111;
    16'b0000010100000001: out_v[143] = 10'b0110001001;
    16'b0000010000000101: out_v[143] = 10'b1001000100;
    16'b0000010100001101: out_v[143] = 10'b0010111101;
    16'b1100010000000001: out_v[143] = 10'b1001000101;
    16'b1100010100001001: out_v[143] = 10'b1101011011;
    16'b0000000000000101: out_v[143] = 10'b1010001101;
    16'b0000000100001001: out_v[143] = 10'b0100111100;
    16'b0100010100001001: out_v[143] = 10'b0010111011;
    16'b0000010100000101: out_v[143] = 10'b1011101010;
    16'b1100000000000101: out_v[143] = 10'b1000001001;
    16'b0100010000000001: out_v[143] = 10'b0001111011;
    16'b1100000100000001: out_v[143] = 10'b1101110011;
    16'b1100000000000001: out_v[143] = 10'b0101100000;
    16'b1000010000000001: out_v[143] = 10'b1101100011;
    16'b0100000100001001: out_v[143] = 10'b0110100011;
    16'b0100010100000001: out_v[143] = 10'b1100011101;
    16'b0000010100001000: out_v[143] = 10'b0110110110;
    16'b0100010000000101: out_v[143] = 10'b0010010111;
    16'b1100010100000101: out_v[143] = 10'b0011111100;
    16'b1000010100000001: out_v[143] = 10'b1011000101;
    16'b1000010000000101: out_v[143] = 10'b0101110010;
    16'b1100010000000100: out_v[143] = 10'b1010111111;
    16'b1100000101001001: out_v[143] = 10'b1011000110;
    16'b1100000100001001: out_v[143] = 10'b0011011101;
    16'b1100000000000100: out_v[143] = 10'b1000001011;
    16'b0000010000000001: out_v[143] = 10'b1001000100;
    16'b1100010100001101: out_v[143] = 10'b1111100010;
    16'b1000010100000101: out_v[143] = 10'b1011001011;
    16'b1000010100001001: out_v[143] = 10'b1011110011;
    16'b0100000100000001: out_v[143] = 10'b0000101111;
    16'b0000000000001001: out_v[143] = 10'b0110000010;
    16'b0000010100000000: out_v[143] = 10'b0111101010;
    16'b0100010100000101: out_v[143] = 10'b1000001011;
    16'b1000000000000101: out_v[143] = 10'b1000111111;
    16'b0100000101001001: out_v[143] = 10'b1101010111;
    16'b0000001000000000: out_v[143] = 10'b0010010000;
    16'b0000001000000001: out_v[143] = 10'b1000110000;
    16'b0000000000000001: out_v[143] = 10'b1110111010;
    16'b0000000000000000: out_v[143] = 10'b0011111000;
    16'b0000001000001001: out_v[143] = 10'b0011001100;
    16'b0000000000001000: out_v[143] = 10'b0111000011;
    16'b0000001100001101: out_v[143] = 10'b1010000000;
    16'b1000001000000000: out_v[143] = 10'b1110010010;
    16'b0000001100001001: out_v[143] = 10'b0001001111;
    16'b0000000100000001: out_v[143] = 10'b0001110011;
    16'b0000000100001101: out_v[143] = 10'b1110110100;
    16'b0010001101001001: out_v[143] = 10'b1010100110;
    16'b0000001101000001: out_v[143] = 10'b0001111010;
    16'b1000010000000100: out_v[143] = 10'b1111011010;
    16'b0010001101000001: out_v[143] = 10'b0110011000;
    16'b0000001100000001: out_v[143] = 10'b1010000101;
    16'b1000011000000100: out_v[143] = 10'b1111010000;
    16'b1000001000000101: out_v[143] = 10'b0011111110;
    16'b1000000100000101: out_v[143] = 10'b0101010100;
    16'b1000000000000100: out_v[143] = 10'b1011100101;
    16'b0000000100000000: out_v[143] = 10'b0011000110;
    16'b1100010001000101: out_v[143] = 10'b1111001011;
    16'b1000000100000001: out_v[143] = 10'b1011001001;
    16'b0000011000000101: out_v[143] = 10'b0000111111;
    16'b1000000000000000: out_v[143] = 10'b1010111001;
    16'b0000001100000000: out_v[143] = 10'b0011000100;
    16'b0010001100000001: out_v[143] = 10'b1010010101;
    16'b1000000001000101: out_v[143] = 10'b0111000110;
    16'b0000000000000100: out_v[143] = 10'b1011101001;
    16'b0010011000000101: out_v[143] = 10'b0010111011;
    16'b1000001101000001: out_v[143] = 10'b0101100010;
    16'b1000011000000101: out_v[143] = 10'b0101100100;
    16'b1000011001000101: out_v[143] = 10'b1010110111;
    16'b1000001000000001: out_v[143] = 10'b0110000011;
    16'b1000010001000101: out_v[143] = 10'b0000011101;
    16'b0000010000000100: out_v[143] = 10'b0100010110;
    16'b0010010000000101: out_v[143] = 10'b1110110110;
    16'b0010001101000000: out_v[143] = 10'b1101100111;
    16'b0000001101000000: out_v[143] = 10'b1111001111;
    16'b1000000000000001: out_v[143] = 10'b0101110000;
    16'b0000011001000101: out_v[143] = 10'b0101101110;
    16'b1000010001000100: out_v[143] = 10'b1111111010;
    16'b1000001100000000: out_v[143] = 10'b1110011010;
    16'b1000001100000001: out_v[143] = 10'b1000110101;
    16'b0000011000000100: out_v[143] = 10'b1010001101;
    16'b1000000001000100: out_v[143] = 10'b1111110101;
    16'b0000001000000101: out_v[143] = 10'b0101101011;
    16'b1000001101000000: out_v[143] = 10'b1101101100;
    16'b0000011100001001: out_v[143] = 10'b0001101100;
    16'b0010010000001001: out_v[143] = 10'b1111001010;
    16'b1000011100000001: out_v[143] = 10'b1111010100;
    16'b0010001100001101: out_v[143] = 10'b0011110010;
    16'b0010010100001001: out_v[143] = 10'b1001001110;
    16'b0010011100001101: out_v[143] = 10'b1010000111;
    16'b1000011100000000: out_v[143] = 10'b0010101000;
    16'b1100011000000101: out_v[143] = 10'b0101001010;
    16'b0000011100001101: out_v[143] = 10'b1100101011;
    16'b0010011000001001: out_v[143] = 10'b1010011010;
    16'b0010011100000101: out_v[143] = 10'b0111110011;
    16'b1000011100001101: out_v[143] = 10'b0111010000;
    16'b1100001000000101: out_v[143] = 10'b0101011010;
    16'b0010001100001001: out_v[143] = 10'b0111010110;
    16'b1010011100001001: out_v[143] = 10'b0100010100;
    16'b1010011100000001: out_v[143] = 10'b1010100011;
    16'b1000011100000101: out_v[143] = 10'b1010011000;
    16'b0000011100000001: out_v[143] = 10'b0100101001;
    16'b0000000100000101: out_v[143] = 10'b1101001110;
    16'b0000011100000101: out_v[143] = 10'b0111001000;
    16'b0010010100001101: out_v[143] = 10'b1010101111;
    16'b0010011100001001: out_v[143] = 10'b0011101100;
    16'b1010011100001101: out_v[143] = 10'b0111111111;
    16'b0010011100000001: out_v[143] = 10'b1100111011;
    16'b0000001100000101: out_v[143] = 10'b0101110010;
    16'b0000001000000100: out_v[143] = 10'b0100111101;
    16'b1000001000000100: out_v[143] = 10'b1111101010;
    16'b1000011100001001: out_v[143] = 10'b0000100110;
    16'b1000001100000101: out_v[143] = 10'b0010100001;
    16'b0000011100001000: out_v[143] = 10'b1011001111;
    16'b1000011000000001: out_v[143] = 10'b0110101111;
    16'b0000011100000000: out_v[143] = 10'b1111110000;
    16'b1000011100000100: out_v[143] = 10'b1111101010;
    16'b0000001100001100: out_v[143] = 10'b0111011010;
    16'b0000001100000100: out_v[143] = 10'b1110111110;
    16'b0000000100000100: out_v[143] = 10'b1010111011;
    16'b0100000000000101: out_v[143] = 10'b1011011000;
    16'b0000001000001000: out_v[143] = 10'b0010010101;
    16'b0000001000001100: out_v[143] = 10'b0000001001;
    16'b0100000000000100: out_v[143] = 10'b1000110010;
    16'b0000001000001101: out_v[143] = 10'b1000100010;
    16'b0000010100001100: out_v[143] = 10'b0101111101;
    16'b0000011000001100: out_v[143] = 10'b0110001011;
    16'b0100000000000000: out_v[143] = 10'b1100100100;
    16'b0000000100001100: out_v[143] = 10'b0111111010;
    16'b0100000000000001: out_v[143] = 10'b0110110010;
    16'b0000011100000100: out_v[143] = 10'b0011111011;
    16'b0000011100001100: out_v[143] = 10'b1000000011;
    16'b0000000000001100: out_v[143] = 10'b1101100001;
    16'b0010010100001100: out_v[143] = 10'b1100000111;
    16'b0010010000000000: out_v[143] = 10'b0001011001;
    16'b0010010000000100: out_v[143] = 10'b0101100111;
    16'b0000010100000100: out_v[143] = 10'b0111001010;
    16'b0000000000001101: out_v[143] = 10'b1101011000;
    16'b0100010100001100: out_v[143] = 10'b0010111111;
    16'b0000010000000000: out_v[143] = 10'b0011010010;
    16'b0010001100001100: out_v[143] = 10'b1111011010;
    16'b0100010000000100: out_v[143] = 10'b0001110111;
    16'b1100000000000000: out_v[143] = 10'b0111000110;
    16'b0100001000000000: out_v[143] = 10'b1000101000;
    16'b0010001001001001: out_v[143] = 10'b1010111010;
    16'b0000010000001001: out_v[143] = 10'b0001100011;
    16'b1000000100001101: out_v[143] = 10'b0100111110;
    16'b0000010000001101: out_v[143] = 10'b0111111101;
    16'b1000010100001101: out_v[143] = 10'b1110011010;
    16'b1100001000000000: out_v[143] = 10'b1000101011;
    16'b0000011000000000: out_v[143] = 10'b1100001111;
    16'b0000011000000001: out_v[143] = 10'b1101001110;
    16'b0100001000000001: out_v[143] = 10'b1011000100;
    16'b0010001000000101: out_v[143] = 10'b1011111011;
    16'b0010001000000001: out_v[143] = 10'b0110000111;
    16'b0010000000000101: out_v[143] = 10'b1111111011;
    16'b0100001100001101: out_v[143] = 10'b1100001111;
    16'b1100001000000001: out_v[143] = 10'b0111010000;
    16'b0100001100001001: out_v[143] = 10'b1101011110;
    16'b0100001000000101: out_v[143] = 10'b1000001101;
    16'b0100000000001001: out_v[143] = 10'b0110111111;
    16'b0100011100001101: out_v[143] = 10'b0110101111;
    16'b0100000100001101: out_v[143] = 10'b1001101010;
    16'b0100010100001101: out_v[143] = 10'b1001100110;
    default: out_v[143] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000000001010: out_v[144] = 10'b1110001011;
    16'b0000010010001000: out_v[144] = 10'b1000010011;
    16'b0000010010011010: out_v[144] = 10'b0010100110;
    16'b0000011010011010: out_v[144] = 10'b1000100001;
    16'b0000010010001010: out_v[144] = 10'b0001101110;
    16'b0000000010001000: out_v[144] = 10'b1100110011;
    16'b0000010000011010: out_v[144] = 10'b1010000011;
    16'b0000011010001000: out_v[144] = 10'b1111100001;
    16'b0000010010011000: out_v[144] = 10'b0010110101;
    16'b0000010000001010: out_v[144] = 10'b0010101111;
    16'b0000010010010010: out_v[144] = 10'b1010011100;
    16'b0000000100001010: out_v[144] = 10'b0111100011;
    16'b0000010010010000: out_v[144] = 10'b1101010011;
    16'b0000000010001010: out_v[144] = 10'b0011111010;
    16'b0000010110011010: out_v[144] = 10'b0100010011;
    16'b0000010100011010: out_v[144] = 10'b1001010100;
    16'b0000000010011010: out_v[144] = 10'b1000100011;
    16'b0000000110001010: out_v[144] = 10'b1011101100;
    16'b0000000000001000: out_v[144] = 10'b1101011011;
    16'b0000001010001000: out_v[144] = 10'b1010100010;
    16'b0000010000010010: out_v[144] = 10'b0001110100;
    16'b0000000010011011: out_v[144] = 10'b0011111111;
    16'b0000001110001000: out_v[144] = 10'b0111011100;
    16'b0000001110000000: out_v[144] = 10'b1000101101;
    16'b0000010000010000: out_v[144] = 10'b0110100001;
    16'b0000000000011010: out_v[144] = 10'b1000100011;
    16'b0000010010000010: out_v[144] = 10'b0100011011;
    16'b0000000000000010: out_v[144] = 10'b0001110111;
    16'b0000000110001000: out_v[144] = 10'b1100111001;
    16'b0000010110001000: out_v[144] = 10'b0100110000;
    16'b0000011010001010: out_v[144] = 10'b0101101000;
    16'b0000010010011011: out_v[144] = 10'b1001100001;
    16'b0000011110011010: out_v[144] = 10'b0110011101;
    16'b0000000010000000: out_v[144] = 10'b0011001111;
    16'b0000011110001000: out_v[144] = 10'b1010101110;
    16'b0000010000000010: out_v[144] = 10'b1101110110;
    16'b0000010000011011: out_v[144] = 10'b0100100011;
    16'b0000010000001000: out_v[144] = 10'b1011011010;
    16'b0000010110001010: out_v[144] = 10'b1010011010;
    16'b0000000110000000: out_v[144] = 10'b1000101010;
    16'b0000000100001000: out_v[144] = 10'b0001011010;
    16'b0000000100000000: out_v[144] = 10'b0010100101;
    16'b0000001010000000: out_v[144] = 10'b1100010011;
    16'b0000000000000000: out_v[144] = 10'b0011011000;
    16'b0000000100001001: out_v[144] = 10'b0100000100;
    16'b0000000100000011: out_v[144] = 10'b0000001100;
    16'b0000010000000000: out_v[144] = 10'b1001100110;
    16'b0000000000000001: out_v[144] = 10'b0010100111;
    16'b0000000100001011: out_v[144] = 10'b0001110101;
    16'b0000010110000000: out_v[144] = 10'b0011011100;
    16'b0000000100000001: out_v[144] = 10'b0110011011;
    16'b0000011110001010: out_v[144] = 10'b0011100101;
    16'b0000001110001010: out_v[144] = 10'b0111010100;
    16'b0000000110000010: out_v[144] = 10'b0011100010;
    16'b0000010100000000: out_v[144] = 10'b1111101010;
    16'b0000011110000000: out_v[144] = 10'b0010111110;
    16'b0000010100001010: out_v[144] = 10'b1010000110;
    16'b0000000100000010: out_v[144] = 10'b0101110100;
    16'b0000000110000001: out_v[144] = 10'b0001101111;
    16'b0000010100001011: out_v[144] = 10'b0001011110;
    16'b0000000110001011: out_v[144] = 10'b1011100011;
    16'b0000001110001011: out_v[144] = 10'b1010001111;
    16'b0000010100001000: out_v[144] = 10'b0000111010;
    16'b0000001110000001: out_v[144] = 10'b0001011001;
    16'b0000010100000001: out_v[144] = 10'b1111000110;
    16'b0000010100000010: out_v[144] = 10'b1011010000;
    16'b0100001110001010: out_v[144] = 10'b0001011111;
    16'b0000000110000011: out_v[144] = 10'b1010111101;
    16'b0000001100000000: out_v[144] = 10'b1011110110;
    16'b0000001110000010: out_v[144] = 10'b0111101110;
    16'b0000001000000000: out_v[144] = 10'b1110111011;
    16'b0100001010000000: out_v[144] = 10'b1000010111;
    16'b0000011010000000: out_v[144] = 10'b0000011111;
    16'b0000001010000010: out_v[144] = 10'b0100011111;
    16'b0000001010001010: out_v[144] = 10'b1011110110;
    16'b0000000010000010: out_v[144] = 10'b0100110111;
    16'b0000010010000000: out_v[144] = 10'b1001011011;
    16'b0000011000000000: out_v[144] = 10'b1110000110;
    16'b0100001010001010: out_v[144] = 10'b1111011011;
    16'b0100011010001010: out_v[144] = 10'b0111011110;
    16'b0000001000001010: out_v[144] = 10'b0111111010;
    16'b0000010000001011: out_v[144] = 10'b0111001010;
    16'b0000010110010010: out_v[144] = 10'b0100010011;
    16'b0000000000010000: out_v[144] = 10'b1111011000;
    16'b0000000000010010: out_v[144] = 10'b1011011010;
    16'b0000000100011010: out_v[144] = 10'b1110111001;
    16'b0000010110010000: out_v[144] = 10'b0011011011;
    16'b0000000010010000: out_v[144] = 10'b1001011011;
    16'b0000000100010000: out_v[144] = 10'b0110100000;
    16'b0000000010010010: out_v[144] = 10'b0110110011;
    16'b0000000110010010: out_v[144] = 10'b0110000001;
    16'b0000000100010010: out_v[144] = 10'b0101111010;
    16'b0000000110010000: out_v[144] = 10'b0000110101;
    16'b0000010110000010: out_v[144] = 10'b0000001101;
    16'b0000010100010010: out_v[144] = 10'b0011111000;
    16'b0000010100010000: out_v[144] = 10'b0111000110;
    16'b0000000110011010: out_v[144] = 10'b1101000010;
    16'b0000001010011010: out_v[144] = 10'b0000101111;
    16'b0000000010001110: out_v[144] = 10'b0011001110;
    16'b0000010100010011: out_v[144] = 10'b1111111011;
    16'b0000000110011000: out_v[144] = 10'b1001101110;
    16'b0000000000011000: out_v[144] = 10'b1011010100;
    default: out_v[144] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1000000000010000: out_v[145] = 10'b0000000011;
    16'b1000000000001000: out_v[145] = 10'b0000001011;
    16'b1000000100001000: out_v[145] = 10'b1000111011;
    16'b1000000100011000: out_v[145] = 10'b0001000001;
    16'b1000000000011000: out_v[145] = 10'b1000100011;
    16'b1100000000000000: out_v[145] = 10'b1011100000;
    16'b1100000000001000: out_v[145] = 10'b0001001001;
    16'b0000000000011000: out_v[145] = 10'b1000110111;
    16'b1100000000010000: out_v[145] = 10'b0010110101;
    16'b0000000000010000: out_v[145] = 10'b0010100011;
    16'b1100000100011000: out_v[145] = 10'b0001110101;
    16'b1100000000111000: out_v[145] = 10'b1111111010;
    16'b1000000100010000: out_v[145] = 10'b0010110011;
    16'b1000000000000000: out_v[145] = 10'b1000110111;
    16'b1100000000011000: out_v[145] = 10'b1011101001;
    16'b1100000100001000: out_v[145] = 10'b0111010011;
    16'b0000000000000000: out_v[145] = 10'b0011100011;
    16'b1000000100000000: out_v[145] = 10'b1111100011;
    16'b0000000100011000: out_v[145] = 10'b0011100111;
    16'b0100000000000000: out_v[145] = 10'b0110010011;
    16'b1000000000111000: out_v[145] = 10'b0110001111;
    16'b0000000000001000: out_v[145] = 10'b1011011101;
    16'b1100100000000000: out_v[145] = 10'b1001111101;
    16'b1100100001000000: out_v[145] = 10'b1001010010;
    16'b0100100001000000: out_v[145] = 10'b0100011100;
    16'b0100100000010000: out_v[145] = 10'b1111001001;
    16'b0100100000000000: out_v[145] = 10'b1100001111;
    16'b1000100001000000: out_v[145] = 10'b0110010111;
    16'b0100100001010000: out_v[145] = 10'b1000101110;
    16'b0000100000000000: out_v[145] = 10'b1000100111;
    16'b0000100000010000: out_v[145] = 10'b1000101100;
    16'b0000100001000000: out_v[145] = 10'b0001010110;
    16'b0000100001010000: out_v[145] = 10'b0010000011;
    16'b1100100001010000: out_v[145] = 10'b1010000111;
    16'b0100000000010000: out_v[145] = 10'b0100111110;
    16'b1100100001110000: out_v[145] = 10'b1001100010;
    16'b1100100001011000: out_v[145] = 10'b1001101100;
    16'b1100100001101000: out_v[145] = 10'b1000110111;
    16'b1100100001100000: out_v[145] = 10'b1110011100;
    16'b0100100101011000: out_v[145] = 10'b0111000000;
    16'b1100100000100000: out_v[145] = 10'b1010101100;
    16'b1100100000101000: out_v[145] = 10'b0110011011;
    16'b0100100001011000: out_v[145] = 10'b0010011001;
    16'b1100100101011000: out_v[145] = 10'b1000101101;
    16'b0100100000011000: out_v[145] = 10'b1111000101;
    16'b0100100001001000: out_v[145] = 10'b0101010110;
    16'b1110100101011000: out_v[145] = 10'b1101010111;
    16'b1100000000101000: out_v[145] = 10'b1110010101;
    16'b0100100001101000: out_v[145] = 10'b0110010010;
    16'b1110100101010000: out_v[145] = 10'b1000111111;
    16'b1100100101000000: out_v[145] = 10'b1011010111;
    16'b1100100001111000: out_v[145] = 10'b1110010111;
    16'b0000100001001000: out_v[145] = 10'b1100011101;
    16'b1100100001001000: out_v[145] = 10'b0010110111;
    16'b1100100101010000: out_v[145] = 10'b1110000100;
    16'b1100100101001000: out_v[145] = 10'b1110011011;
    16'b1100100000010000: out_v[145] = 10'b0101011111;
    16'b1100100000110000: out_v[145] = 10'b1011100010;
    16'b1100100000011000: out_v[145] = 10'b1011010101;
    16'b1100100000111000: out_v[145] = 10'b1001010010;
    16'b1100000000100000: out_v[145] = 10'b1100011011;
    16'b0100100001100000: out_v[145] = 10'b1111100101;
    16'b1100100100011000: out_v[145] = 10'b0111111010;
    16'b1100100000001000: out_v[145] = 10'b0111000110;
    16'b1000100001010000: out_v[145] = 10'b0110110001;
    16'b1100100100010000: out_v[145] = 10'b0110101110;
    16'b0000100001011000: out_v[145] = 10'b0100011111;
    16'b0100100000001000: out_v[145] = 10'b1011100110;
    16'b0000000101011000: out_v[145] = 10'b1001100111;
    16'b1000100000000000: out_v[145] = 10'b1101010000;
    16'b1000000001011000: out_v[145] = 10'b0111101110;
    16'b1000000001001000: out_v[145] = 10'b0101000100;
    16'b1000100001011000: out_v[145] = 10'b0000001110;
    16'b1000000001000000: out_v[145] = 10'b1011001100;
    16'b0000000001011000: out_v[145] = 10'b1000100111;
    16'b0000100101011000: out_v[145] = 10'b1001001010;
    16'b1000000101011000: out_v[145] = 10'b0001001111;
    16'b1000000001010000: out_v[145] = 10'b1111110011;
    16'b0000100100011000: out_v[145] = 10'b1001001001;
    16'b1100000001000000: out_v[145] = 10'b1101101100;
    16'b1000100101011000: out_v[145] = 10'b0000111001;
    16'b0000100000011000: out_v[145] = 10'b1000111100;
    16'b1000100101010000: out_v[145] = 10'b1100011111;
    16'b1100000001010000: out_v[145] = 10'b0100101100;
    16'b0000000001000000: out_v[145] = 10'b1101010010;
    16'b1000100001001000: out_v[145] = 10'b1111001011;
    16'b1100000001011000: out_v[145] = 10'b1010111010;
    16'b1100000001101000: out_v[145] = 10'b1010011111;
    16'b0000000001010000: out_v[145] = 10'b0110111110;
    16'b0000100000001000: out_v[145] = 10'b0000111110;
    16'b1000100000011000: out_v[145] = 10'b0111100100;
    16'b1000000001101000: out_v[145] = 10'b1010101101;
    16'b1100000001001000: out_v[145] = 10'b1100110011;
    16'b0000100101010000: out_v[145] = 10'b1001101011;
    16'b0000000001001000: out_v[145] = 10'b0001111100;
    16'b1000100000010000: out_v[145] = 10'b1010110000;
    16'b1000100000001000: out_v[145] = 10'b1001101111;
    16'b1000000101001000: out_v[145] = 10'b1111100000;
    16'b0000100101001000: out_v[145] = 10'b0100011111;
    16'b0000100101000000: out_v[145] = 10'b0010110101;
    16'b0000000101000000: out_v[145] = 10'b0101010011;
    16'b0000100100001000: out_v[145] = 10'b0001111010;
    16'b0000100100000000: out_v[145] = 10'b0011010101;
    16'b0100100101000000: out_v[145] = 10'b0011110011;
    16'b1000000101010000: out_v[145] = 10'b0100000110;
    16'b1000100100011000: out_v[145] = 10'b0110111011;
    16'b1100000001111000: out_v[145] = 10'b1110100111;
    16'b0100100101001001: out_v[145] = 10'b1111101111;
    16'b1100100101001001: out_v[145] = 10'b1110101110;
    16'b1000100001111000: out_v[145] = 10'b1101010110;
    16'b0100100001111000: out_v[145] = 10'b0100100110;
    16'b1000000001111000: out_v[145] = 10'b0111000011;
    16'b0100100000111000: out_v[145] = 10'b0011100111;
    16'b0100100000110000: out_v[145] = 10'b1011111001;
    16'b0100100001110000: out_v[145] = 10'b1001001110;
    16'b1100100101111000: out_v[145] = 10'b1000110010;
    16'b1000100000111000: out_v[145] = 10'b1101001110;
    16'b0100100101001000: out_v[145] = 10'b1111101001;
    16'b1100100100000000: out_v[145] = 10'b0110101111;
    16'b0000000100001000: out_v[145] = 10'b1010010000;
    16'b0000000100010000: out_v[145] = 10'b1101110011;
    16'b0100100101010000: out_v[145] = 10'b1111001111;
    16'b1100000100010000: out_v[145] = 10'b0011000110;
    16'b0000000100000000: out_v[145] = 10'b1110000010;
    16'b1100000100000000: out_v[145] = 10'b0011111011;
    16'b0000000101010000: out_v[145] = 10'b0100001111;
    16'b0100000100010000: out_v[145] = 10'b0100110110;
    16'b0001000100000000: out_v[145] = 10'b1010011001;
    16'b0100100100000000: out_v[145] = 10'b0101011010;
    16'b0100000100000000: out_v[145] = 10'b0000111111;
    16'b0001001100000000: out_v[145] = 10'b0101011011;
    16'b1000100101000000: out_v[145] = 10'b0110001010;
    16'b1000100101001000: out_v[145] = 10'b1111011010;
    16'b0100000100011000: out_v[145] = 10'b1000100111;
    16'b0000100100010000: out_v[145] = 10'b1001011110;
    default: out_v[145] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001000010000000: out_v[146] = 10'b0000011101;
    16'b0001000010100000: out_v[146] = 10'b0110100001;
    16'b0000000000000000: out_v[146] = 10'b1011100110;
    16'b0001000000000000: out_v[146] = 10'b0101001110;
    16'b0000000010000000: out_v[146] = 10'b1100000111;
    16'b0001000000100000: out_v[146] = 10'b0000011001;
    16'b0000000110000000: out_v[146] = 10'b0110110111;
    16'b0001000110000000: out_v[146] = 10'b1010100000;
    16'b0000000010100000: out_v[146] = 10'b1100100001;
    16'b0000000100000000: out_v[146] = 10'b1000111101;
    16'b0001000000010000: out_v[146] = 10'b0001010100;
    16'b0001000010000001: out_v[146] = 10'b0100001110;
    16'b0001000010010000: out_v[146] = 10'b0000011111;
    16'b0000000000010000: out_v[146] = 10'b1110000111;
    16'b0000000010010000: out_v[146] = 10'b1010010110;
    16'b0000000000100000: out_v[146] = 10'b0010011110;
    16'b0000000010000001: out_v[146] = 10'b0010101110;
    16'b0001000100010000: out_v[146] = 10'b0111001010;
    16'b0001000100000000: out_v[146] = 10'b1111100000;
    16'b0001000010000011: out_v[146] = 10'b0111001001;
    16'b0001000110010000: out_v[146] = 10'b1011111011;
    16'b0001000100100000: out_v[146] = 10'b0110010101;
    16'b0000000110100000: out_v[146] = 10'b0000110110;
    16'b0001000110100000: out_v[146] = 10'b1111100011;
    16'b0001000000000100: out_v[146] = 10'b1101110110;
    16'b0001000010000100: out_v[146] = 10'b0001010010;
    16'b0000000000000100: out_v[146] = 10'b1010100000;
    16'b0000000010000100: out_v[146] = 10'b1101011001;
    16'b0100000010100000: out_v[146] = 10'b1001111101;
    16'b0100000010000000: out_v[146] = 10'b1111001000;
    16'b0100000000000000: out_v[146] = 10'b1111100110;
    default: out_v[146] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001001101010001: out_v[147] = 10'b1110100011;
    16'b0001000101010000: out_v[147] = 10'b1011010001;
    16'b0001000101000000: out_v[147] = 10'b1011110010;
    16'b0000000101010001: out_v[147] = 10'b0011110000;
    16'b0101000101010000: out_v[147] = 10'b0111100111;
    16'b0000000101000000: out_v[147] = 10'b0011100111;
    16'b0001000100000000: out_v[147] = 10'b0010101011;
    16'b0000000000000000: out_v[147] = 10'b0001011110;
    16'b0000000001010001: out_v[147] = 10'b0001010101;
    16'b0101000101000000: out_v[147] = 10'b1001110010;
    16'b0101001101010000: out_v[147] = 10'b0111110011;
    16'b0001000101010001: out_v[147] = 10'b0010101011;
    16'b0000000101000001: out_v[147] = 10'b1010110010;
    16'b0100000101000001: out_v[147] = 10'b0000011101;
    16'b0001000101000001: out_v[147] = 10'b1011001100;
    16'b0000000001000001: out_v[147] = 10'b1110100001;
    16'b0001000100000001: out_v[147] = 10'b1100011111;
    16'b0000000100000000: out_v[147] = 10'b0110001011;
    16'b0000000101010000: out_v[147] = 10'b1101100100;
    16'b0000000100000001: out_v[147] = 10'b0010011111;
    16'b0000000001010000: out_v[147] = 10'b0000001111;
    16'b0100000101000000: out_v[147] = 10'b1001011001;
    16'b0001000000000000: out_v[147] = 10'b1001101110;
    16'b0001000001000000: out_v[147] = 10'b0011110101;
    16'b0100000101010001: out_v[147] = 10'b1010110001;
    16'b0101000101000001: out_v[147] = 10'b1111001100;
    16'b0101001100000001: out_v[147] = 10'b0101000011;
    16'b0101000101010001: out_v[147] = 10'b0001101100;
    16'b0001001101010000: out_v[147] = 10'b1010000110;
    16'b0001000100010000: out_v[147] = 10'b0100100101;
    16'b0100001001000000: out_v[147] = 10'b1011100010;
    16'b0100000001010000: out_v[147] = 10'b0101011000;
    16'b0000000000010000: out_v[147] = 10'b1100001111;
    16'b0000001001010000: out_v[147] = 10'b0110111000;
    16'b0000000100010000: out_v[147] = 10'b0110001111;
    16'b0000001100010000: out_v[147] = 10'b0111010001;
    16'b0100000100000001: out_v[147] = 10'b1001010101;
    16'b0000001001000000: out_v[147] = 10'b1011011110;
    16'b0100000100010000: out_v[147] = 10'b1010100110;
    16'b0100001001010000: out_v[147] = 10'b0100110011;
    16'b0000001101010000: out_v[147] = 10'b0001011110;
    16'b0100000000010000: out_v[147] = 10'b1001001110;
    16'b0100001000000000: out_v[147] = 10'b0000101111;
    16'b0100000100000000: out_v[147] = 10'b1111000001;
    16'b0100000001000000: out_v[147] = 10'b1101000010;
    16'b0100000000000000: out_v[147] = 10'b0101111000;
    16'b0000001000010000: out_v[147] = 10'b1001110011;
    16'b0100001101010000: out_v[147] = 10'b0000011110;
    16'b0100001000010000: out_v[147] = 10'b0010111111;
    16'b0100001100010000: out_v[147] = 10'b0010001101;
    16'b0000000001000000: out_v[147] = 10'b1111100001;
    16'b0100001100000001: out_v[147] = 10'b0110100000;
    16'b0100001101000001: out_v[147] = 10'b1101100100;
    16'b0000001000000000: out_v[147] = 10'b0010110101;
    16'b0100001101010001: out_v[147] = 10'b1001100100;
    16'b0100001001010001: out_v[147] = 10'b1011100100;
    16'b0000001100000000: out_v[147] = 10'b0010110101;
    16'b0100001001000001: out_v[147] = 10'b1111100110;
    16'b0100000001010001: out_v[147] = 10'b1010001101;
    16'b0100000001000001: out_v[147] = 10'b1111101000;
    16'b0000001100010001: out_v[147] = 10'b1110001001;
    16'b0100001000010001: out_v[147] = 10'b1111010100;
    16'b0000001000010001: out_v[147] = 10'b1011000100;
    16'b0100001101010011: out_v[147] = 10'b0111010111;
    16'b0000001101010001: out_v[147] = 10'b1111010100;
    16'b0100001100000000: out_v[147] = 10'b1000000110;
    16'b0100000101010000: out_v[147] = 10'b0100011101;
    16'b0000001101000001: out_v[147] = 10'b1101100110;
    16'b0100001100010001: out_v[147] = 10'b0100010001;
    16'b0100000000010001: out_v[147] = 10'b0011101001;
    16'b0001001100000001: out_v[147] = 10'b1011101011;
    16'b0100001101000000: out_v[147] = 10'b0110000001;
    16'b0000001001010001: out_v[147] = 10'b0111111000;
    16'b0000001100000001: out_v[147] = 10'b0110101111;
    16'b0000001001000001: out_v[147] = 10'b1110011110;
    16'b0101000001010001: out_v[147] = 10'b1010001000;
    16'b0101000100000001: out_v[147] = 10'b0010011100;
    16'b0001000001000001: out_v[147] = 10'b1010110000;
    16'b0101000100000000: out_v[147] = 10'b1011000011;
    16'b0101000001010000: out_v[147] = 10'b0110001101;
    16'b0101000001000001: out_v[147] = 10'b1100000110;
    16'b0001000001010001: out_v[147] = 10'b1000001110;
    16'b0111000101000001: out_v[147] = 10'b0001011111;
    16'b0101001000010000: out_v[147] = 10'b0100111110;
    16'b0101000000000000: out_v[147] = 10'b0010010001;
    16'b0001001100000000: out_v[147] = 10'b1100011000;
    16'b0110000010000000: out_v[147] = 10'b0000111011;
    16'b0100000010000000: out_v[147] = 10'b0000100111;
    16'b0101000001000000: out_v[147] = 10'b1010110111;
    16'b0101001000000000: out_v[147] = 10'b1111110100;
    16'b0110000000010000: out_v[147] = 10'b0011111111;
    16'b0110001000000000: out_v[147] = 10'b0111111111;
    16'b0101000010000000: out_v[147] = 10'b0011111100;
    16'b0111000000000000: out_v[147] = 10'b0000110011;
    16'b0110000000000000: out_v[147] = 10'b1101001101;
    16'b0010000000000000: out_v[147] = 10'b1111010000;
    16'b0101001001000000: out_v[147] = 10'b1100010000;
    16'b0001001000000000: out_v[147] = 10'b1101000001;
    16'b0010001000000000: out_v[147] = 10'b1001010111;
    16'b0101001100000000: out_v[147] = 10'b1100110101;
    16'b0101001101000000: out_v[147] = 10'b0100110111;
    16'b0101000000000001: out_v[147] = 10'b1101001000;
    16'b0101000000010000: out_v[147] = 10'b0001111101;
    16'b0101000100010000: out_v[147] = 10'b1101000000;
    16'b0101001100010000: out_v[147] = 10'b1011001100;
    16'b0111001000000000: out_v[147] = 10'b1011110011;
    16'b0001001001000000: out_v[147] = 10'b1001011000;
    16'b0001001101000000: out_v[147] = 10'b0110110011;
    16'b0001000100010001: out_v[147] = 10'b0110101101;
    16'b0101000100010001: out_v[147] = 10'b1110100010;
    16'b0001000100010010: out_v[147] = 10'b1110001010;
    16'b0101001100010001: out_v[147] = 10'b1011010011;
    16'b0001000101010010: out_v[147] = 10'b1111001010;
    16'b0100000000000001: out_v[147] = 10'b1111001000;
    16'b0001001100010000: out_v[147] = 10'b1011011000;
    16'b0101001101010010: out_v[147] = 10'b0011111110;
    16'b0100001000000001: out_v[147] = 10'b1101010100;
    16'b0101001000000001: out_v[147] = 10'b0011100110;
    16'b0001001100010010: out_v[147] = 10'b0100111111;
    16'b0001001101010010: out_v[147] = 10'b1101011101;
    16'b0101000100010010: out_v[147] = 10'b1101011110;
    16'b0001001100010001: out_v[147] = 10'b1011010101;
    16'b0000000000000001: out_v[147] = 10'b0110011001;
    16'b0101001100010010: out_v[147] = 10'b0011000110;
    16'b0000001000000001: out_v[147] = 10'b0110110000;
    16'b0001001000000001: out_v[147] = 10'b1100010010;
    16'b0110010010000000: out_v[147] = 10'b1110000101;
    16'b0100000110000000: out_v[147] = 10'b1011100001;
    16'b0100010110000000: out_v[147] = 10'b1010100010;
    16'b0100010010000000: out_v[147] = 10'b0111011101;
    16'b0100001110000000: out_v[147] = 10'b1001101011;
    16'b0000000010000000: out_v[147] = 10'b0110011110;
    16'b0110010110000000: out_v[147] = 10'b0110001111;
    16'b0110000110000000: out_v[147] = 10'b0101011110;
    16'b0101001001010001: out_v[147] = 10'b1100101010;
    16'b0101001101010001: out_v[147] = 10'b0111011011;
    16'b0101001000010001: out_v[147] = 10'b1011000110;
    16'b0101001101000001: out_v[147] = 10'b0111100000;
    16'b0111001100000001: out_v[147] = 10'b1111101001;
    16'b0101000000010001: out_v[147] = 10'b1110100010;
    16'b0110001100000000: out_v[147] = 10'b1010011000;
    16'b0110001110000000: out_v[147] = 10'b1101001010;
    16'b0101000110000000: out_v[147] = 10'b1101101010;
    16'b0111001110000000: out_v[147] = 10'b1111001011;
    16'b0111000110000000: out_v[147] = 10'b1101100011;
    16'b0100011110000000: out_v[147] = 10'b1101101011;
    16'b0110000100000000: out_v[147] = 10'b1111010101;
    16'b0101001110000000: out_v[147] = 10'b0110101100;
    default: out_v[147] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000101000000100: out_v[148] = 10'b0000000111;
    16'b0000101000010000: out_v[148] = 10'b1111011100;
    16'b0000101000011000: out_v[148] = 10'b0101010000;
    16'b1100101000000000: out_v[148] = 10'b0101100111;
    16'b0000101000000000: out_v[148] = 10'b1010100101;
    16'b0100101000010000: out_v[148] = 10'b1001011000;
    16'b0000100000000000: out_v[148] = 10'b1010000011;
    16'b0000001000011000: out_v[148] = 10'b1110001011;
    16'b0000101000001000: out_v[148] = 10'b1111100000;
    16'b1000101000010000: out_v[148] = 10'b0000011011;
    16'b0100001000010000: out_v[148] = 10'b0110011110;
    16'b1000001000011000: out_v[148] = 10'b0111010011;
    16'b0000001000010000: out_v[148] = 10'b1111100100;
    16'b0000000000010000: out_v[148] = 10'b0100110010;
    16'b0100101000000000: out_v[148] = 10'b0100110101;
    16'b0000100000000100: out_v[148] = 10'b1110001001;
    16'b1000101000000000: out_v[148] = 10'b1010111000;
    16'b1000101000011000: out_v[148] = 10'b1001111011;
    16'b0000001000000000: out_v[148] = 10'b0111001100;
    16'b1100001000010000: out_v[148] = 10'b1100100101;
    16'b1100101000010000: out_v[148] = 10'b0111101111;
    16'b0000001000011100: out_v[148] = 10'b0100101011;
    16'b1000001000010000: out_v[148] = 10'b1100110100;
    16'b0000101000011100: out_v[148] = 10'b1011001001;
    16'b0000001000000100: out_v[148] = 10'b1101110101;
    16'b0000101000001100: out_v[148] = 10'b0011100110;
    16'b0000000000000000: out_v[148] = 10'b1001001110;
    16'b0000101000010100: out_v[148] = 10'b1000101101;
    16'b1000101000001000: out_v[148] = 10'b1111100111;
    16'b0000000000000100: out_v[148] = 10'b1110111010;
    16'b0000100000010000: out_v[148] = 10'b0110011010;
    16'b1000100000010000: out_v[148] = 10'b1101010110;
    16'b0100100000000000: out_v[148] = 10'b1110110111;
    16'b1100100000000000: out_v[148] = 10'b1101010110;
    16'b1100100000110000: out_v[148] = 10'b0101110110;
    16'b1000100000000000: out_v[148] = 10'b1100011100;
    16'b1100100000010000: out_v[148] = 10'b1111100101;
    16'b1100101000110000: out_v[148] = 10'b1101011000;
    16'b1100000000010000: out_v[148] = 10'b1001101111;
    16'b1000000000000000: out_v[148] = 10'b0100111100;
    16'b1000001000000000: out_v[148] = 10'b0101100011;
    16'b1100101000100000: out_v[148] = 10'b0110001111;
    16'b0000101000010010: out_v[148] = 10'b0001011011;
    16'b1000100000000100: out_v[148] = 10'b0111010111;
    16'b1000101000000100: out_v[148] = 10'b1011111011;
    16'b0000100000010100: out_v[148] = 10'b0101010000;
    16'b0000000000010100: out_v[148] = 10'b1110100010;
    16'b0000001000010100: out_v[148] = 10'b1000100011;
    16'b0000000000001000: out_v[148] = 10'b0001100111;
    16'b0000100000001000: out_v[148] = 10'b0100110101;
    16'b0001000000000000: out_v[148] = 10'b1101001111;
    16'b0000001000001000: out_v[148] = 10'b1101111010;
    16'b0000010000000000: out_v[148] = 10'b0011000011;
    16'b0010101000000000: out_v[148] = 10'b1101011101;
    16'b0010100000000000: out_v[148] = 10'b1010101011;
    default: out_v[148] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000010000001000: out_v[149] = 10'b1000001011;
    16'b0100010000001000: out_v[149] = 10'b0110100011;
    16'b1001010010001000: out_v[149] = 10'b0111100110;
    16'b0000010000001010: out_v[149] = 10'b1011101010;
    16'b1001010010000000: out_v[149] = 10'b0111010010;
    16'b0101000010001000: out_v[149] = 10'b0001011110;
    16'b1001000010000000: out_v[149] = 10'b1010100010;
    16'b0000000000001000: out_v[149] = 10'b1010100001;
    16'b0000010000001011: out_v[149] = 10'b1101111001;
    16'b1001010001001000: out_v[149] = 10'b1101000111;
    16'b0000010000000000: out_v[149] = 10'b0110011011;
    16'b0000010001001000: out_v[149] = 10'b0000010111;
    16'b0001010010001000: out_v[149] = 10'b1011001110;
    16'b0100000000001000: out_v[149] = 10'b0010101010;
    16'b1001010011001000: out_v[149] = 10'b0100010101;
    16'b1001000010001000: out_v[149] = 10'b0001011101;
    16'b0001010000001000: out_v[149] = 10'b1100001001;
    16'b1001010011000000: out_v[149] = 10'b0100011011;
    16'b0100010000001010: out_v[149] = 10'b1001010100;
    16'b0000010000001001: out_v[149] = 10'b1011010111;
    16'b1101000010001000: out_v[149] = 10'b1010010111;
    16'b1000000011001000: out_v[149] = 10'b1010101011;
    16'b0100010000001001: out_v[149] = 10'b1010111010;
    16'b0101010010001000: out_v[149] = 10'b0111010011;
    16'b0001000000001000: out_v[149] = 10'b0010011011;
    16'b0000000000000000: out_v[149] = 10'b0011100001;
    16'b1001000011001000: out_v[149] = 10'b0000110101;
    16'b1101010010001000: out_v[149] = 10'b0110110111;
    16'b0001000010001000: out_v[149] = 10'b1011011110;
    16'b0000000000001010: out_v[149] = 10'b1011101110;
    16'b0000010000000011: out_v[149] = 10'b0010110101;
    16'b0100010000001011: out_v[149] = 10'b1100011110;
    16'b1001010010001010: out_v[149] = 10'b1111001000;
    16'b1001010010001001: out_v[149] = 10'b1011010111;
    16'b1001010000001000: out_v[149] = 10'b1101011010;
    16'b0100010000000011: out_v[149] = 10'b1110011011;
    16'b0001010001001000: out_v[149] = 10'b1100010011;
    16'b0001000010000000: out_v[149] = 10'b0110011001;
    16'b0001010010001010: out_v[149] = 10'b1001100011;
    16'b1000010011001000: out_v[149] = 10'b0101100011;
    16'b0100000000000001: out_v[149] = 10'b1101100111;
    16'b0000000000000011: out_v[149] = 10'b1000100010;
    16'b0000000000000001: out_v[149] = 10'b0100100110;
    16'b0000000000001011: out_v[149] = 10'b1000101011;
    16'b0000000000001001: out_v[149] = 10'b0111001000;
    16'b0100000000000011: out_v[149] = 10'b0111011010;
    16'b0000000001000011: out_v[149] = 10'b0110000101;
    16'b0000000001101011: out_v[149] = 10'b1001111001;
    16'b0000010001001010: out_v[149] = 10'b0001110111;
    16'b0000000001000010: out_v[149] = 10'b0000011010;
    16'b0000000001001010: out_v[149] = 10'b0111010010;
    16'b0000000001001001: out_v[149] = 10'b0001111010;
    16'b1000000001001011: out_v[149] = 10'b0101011101;
    16'b0000000000000010: out_v[149] = 10'b0010110000;
    16'b1000000001001010: out_v[149] = 10'b1100101011;
    16'b0100010000000010: out_v[149] = 10'b1011110100;
    16'b0000000001101001: out_v[149] = 10'b1101000001;
    16'b0000010001101010: out_v[149] = 10'b1100111111;
    16'b0000000001001011: out_v[149] = 10'b0011011001;
    16'b0000010000000010: out_v[149] = 10'b1100111000;
    16'b1000010001001010: out_v[149] = 10'b0011110100;
    16'b0000000001001000: out_v[149] = 10'b0001011110;
    16'b0000010001000010: out_v[149] = 10'b1001001010;
    16'b0000000001101010: out_v[149] = 10'b0111111011;
    16'b0000000001000001: out_v[149] = 10'b1100001000;
    16'b0100000000001010: out_v[149] = 10'b1001100110;
    16'b1000000001001001: out_v[149] = 10'b0001001111;
    16'b0000010001001001: out_v[149] = 10'b0111011000;
    16'b0000000001000000: out_v[149] = 10'b0001011110;
    16'b1000000001000001: out_v[149] = 10'b0000011101;
    16'b0100000000001011: out_v[149] = 10'b0111101000;
    16'b0000000011001001: out_v[149] = 10'b0111001111;
    16'b0000010001001011: out_v[149] = 10'b0110010111;
    16'b0000010001000001: out_v[149] = 10'b0101001010;
    16'b0100000001001001: out_v[149] = 10'b0010111011;
    16'b0100000000001001: out_v[149] = 10'b1100000111;
    16'b1000010001001001: out_v[149] = 10'b0001111100;
    16'b1000000000001001: out_v[149] = 10'b0011111110;
    16'b0001000000001010: out_v[149] = 10'b1011001010;
    16'b1001000011000010: out_v[149] = 10'b0111001011;
    16'b0000010010000010: out_v[149] = 10'b1100000100;
    16'b1001010011000010: out_v[149] = 10'b0011111110;
    16'b1001000010000010: out_v[149] = 10'b1101111111;
    16'b0100000000000010: out_v[149] = 10'b0000111000;
    16'b1001010001000010: out_v[149] = 10'b0001010110;
    16'b0100010010000010: out_v[149] = 10'b1111011011;
    16'b0101010010000010: out_v[149] = 10'b1111111111;
    16'b1001010010000010: out_v[149] = 10'b1101001011;
    16'b0001000000000010: out_v[149] = 10'b1011011110;
    16'b0100000010000010: out_v[149] = 10'b1111111101;
    16'b1001000000001010: out_v[149] = 10'b0111000111;
    16'b1001000001000010: out_v[149] = 10'b0101110010;
    16'b0001010000000010: out_v[149] = 10'b1101000011;
    16'b0001010010000010: out_v[149] = 10'b1101001111;
    16'b1101010010000010: out_v[149] = 10'b0011110001;
    16'b0101000010000010: out_v[149] = 10'b0011001111;
    16'b1001000010001010: out_v[149] = 10'b0111000110;
    16'b0000000010001010: out_v[149] = 10'b0111111110;
    16'b0000000010000010: out_v[149] = 10'b0111001101;
    16'b1101010011000010: out_v[149] = 10'b1010011010;
    16'b1001000000000010: out_v[149] = 10'b1001001010;
    16'b0001000001000010: out_v[149] = 10'b1111000010;
    16'b1101000010000010: out_v[149] = 10'b0111011110;
    16'b0001000010000010: out_v[149] = 10'b0110010001;
    16'b1101000010001001: out_v[149] = 10'b0111101011;
    16'b0001000000001001: out_v[149] = 10'b0110011100;
    16'b0101000000001001: out_v[149] = 10'b1110001110;
    16'b1001000001001001: out_v[149] = 10'b1111110111;
    16'b1001000011001001: out_v[149] = 10'b0010111111;
    16'b0001000001001001: out_v[149] = 10'b1001111111;
    16'b1001010001001001: out_v[149] = 10'b0111010100;
    16'b1001010011001001: out_v[149] = 10'b1110110100;
    16'b1001000000001001: out_v[149] = 10'b0100110010;
    16'b1101000001001001: out_v[149] = 10'b1010110111;
    16'b1101000011001001: out_v[149] = 10'b0000111101;
    16'b1101000000001001: out_v[149] = 10'b0010011111;
    16'b0000010000000001: out_v[149] = 10'b0011100010;
    16'b1001010011000011: out_v[149] = 10'b0101010110;
    16'b0001010000000000: out_v[149] = 10'b0111111110;
    16'b1001010001000001: out_v[149] = 10'b0101110100;
    16'b0001010001000010: out_v[149] = 10'b0000111101;
    16'b1001010011000001: out_v[149] = 10'b0001001011;
    16'b1011010000000010: out_v[149] = 10'b1010111101;
    16'b1001010000000010: out_v[149] = 10'b0001111111;
    16'b1000010000000010: out_v[149] = 10'b0011110000;
    16'b1000000000000010: out_v[149] = 10'b0111011010;
    16'b1010010000000000: out_v[149] = 10'b1110110111;
    16'b1000000000000011: out_v[149] = 10'b1111000011;
    16'b1010000000000010: out_v[149] = 10'b0101100111;
    16'b1011010010000011: out_v[149] = 10'b0011111110;
    16'b1010010000000010: out_v[149] = 10'b1110101001;
    16'b1011010000000000: out_v[149] = 10'b0101110101;
    16'b1001010010000011: out_v[149] = 10'b1110101001;
    16'b1001010000000000: out_v[149] = 10'b0010011111;
    16'b1000000000000000: out_v[149] = 10'b1110100110;
    16'b1011000000000010: out_v[149] = 10'b1011101011;
    16'b1001000000000011: out_v[149] = 10'b0010001001;
    16'b1000000000001010: out_v[149] = 10'b0111011010;
    16'b1001000000000000: out_v[149] = 10'b1011110111;
    16'b1011010010000010: out_v[149] = 10'b0001111110;
    16'b1001010000000011: out_v[149] = 10'b0101001010;
    16'b1011010000000011: out_v[149] = 10'b0111000111;
    16'b1001010001001010: out_v[149] = 10'b1101001010;
    16'b0001000000001011: out_v[149] = 10'b1110001011;
    16'b1001010001001011: out_v[149] = 10'b1101001011;
    16'b1001000001001010: out_v[149] = 10'b0110111010;
    16'b1001000001001011: out_v[149] = 10'b1000100111;
    16'b1001010000001010: out_v[149] = 10'b1111100011;
    16'b1001000000001011: out_v[149] = 10'b0100011001;
    16'b0001000000000011: out_v[149] = 10'b1110000101;
    16'b0001010000001011: out_v[149] = 10'b0101011111;
    16'b1001010010001011: out_v[149] = 10'b1001011011;
    16'b0001010000000011: out_v[149] = 10'b0001011010;
    16'b0001010000001010: out_v[149] = 10'b1101000010;
    16'b1001000010000001: out_v[149] = 10'b1100101100;
    16'b0001000000000001: out_v[149] = 10'b1101000101;
    16'b1001000010001011: out_v[149] = 10'b1101010011;
    16'b0001000000000000: out_v[149] = 10'b1000101111;
    16'b1001000010000011: out_v[149] = 10'b1001100100;
    default: out_v[149] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000110010000: out_v[150] = 10'b1000000111;
    16'b0000100100010010: out_v[150] = 10'b1001100011;
    16'b0000100000010010: out_v[150] = 10'b0010100010;
    16'b0000000100010010: out_v[150] = 10'b0011101100;
    16'b0000000100010000: out_v[150] = 10'b1100100001;
    16'b0000000000110010: out_v[150] = 10'b0011110001;
    16'b0000100000010000: out_v[150] = 10'b0110011000;
    16'b0000000000000010: out_v[150] = 10'b0010000110;
    16'b0000100100000010: out_v[150] = 10'b0100000001;
    16'b0000100100100010: out_v[150] = 10'b0000011111;
    16'b0000000100000000: out_v[150] = 10'b0011001000;
    16'b0000000110110010: out_v[150] = 10'b1100110001;
    16'b0000000100110010: out_v[150] = 10'b0011111100;
    16'b0000000000010000: out_v[150] = 10'b0101111011;
    16'b0000100000000010: out_v[150] = 10'b1111000011;
    16'b0000000110010010: out_v[150] = 10'b0111000001;
    16'b0000000010110010: out_v[150] = 10'b0000111001;
    16'b0000000000010010: out_v[150] = 10'b0011100111;
    16'b0000100100010000: out_v[150] = 10'b1100001001;
    16'b0000100110100010: out_v[150] = 10'b1100010111;
    16'b0000100110110010: out_v[150] = 10'b0000010111;
    16'b0000000110100010: out_v[150] = 10'b0010101001;
    16'b0000000100000010: out_v[150] = 10'b0110010011;
    16'b0000000100100010: out_v[150] = 10'b0101001010;
    16'b0000100100110010: out_v[150] = 10'b1011101110;
    16'b0000000000000000: out_v[150] = 10'b0111011000;
    16'b0000000000100010: out_v[150] = 10'b0001001010;
    16'b0000000010000000: out_v[150] = 10'b1001011110;
    16'b0000000000100001: out_v[150] = 10'b1110100100;
    16'b0000000100010001: out_v[150] = 10'b1100111010;
    16'b0000000000100000: out_v[150] = 10'b1011000111;
    16'b0000000100100000: out_v[150] = 10'b0010100111;
    16'b0000000010100000: out_v[150] = 10'b1101001010;
    16'b0000000100100001: out_v[150] = 10'b0110000101;
    16'b0000000110000000: out_v[150] = 10'b0011001101;
    16'b0000000110100000: out_v[150] = 10'b1001101000;
    16'b0000100100110000: out_v[150] = 10'b1100000110;
    16'b0000000100110000: out_v[150] = 10'b0010010101;
    16'b0000000000110000: out_v[150] = 10'b1000010111;
    16'b0000000100110001: out_v[150] = 10'b0000111101;
    16'b0000000000000001: out_v[150] = 10'b1010011101;
    16'b0000000100000001: out_v[150] = 10'b0110011001;
    16'b0000000110110000: out_v[150] = 10'b0110010001;
    16'b0000000010100010: out_v[150] = 10'b0100001000;
    16'b0000000010010000: out_v[150] = 10'b1000010100;
    16'b0000000010000010: out_v[150] = 10'b0111100110;
    16'b0000000110000010: out_v[150] = 10'b1001110010;
    16'b0000000010010010: out_v[150] = 10'b0110110100;
    16'b0000100000000000: out_v[150] = 10'b0000100000;
    16'b0000100100000000: out_v[150] = 10'b0010100110;
    16'b0000100010000000: out_v[150] = 10'b0001100110;
    16'b0000000000110011: out_v[150] = 10'b1011100010;
    16'b0000000000010011: out_v[150] = 10'b1011000010;
    16'b0000000000100011: out_v[150] = 10'b1001001010;
    16'b0000000000010001: out_v[150] = 10'b1001101000;
    16'b0000000000000011: out_v[150] = 10'b1011100110;
    16'b0001010010010000: out_v[150] = 10'b0101110110;
    16'b0000100110010000: out_v[150] = 10'b0110011001;
    16'b0001000010000000: out_v[150] = 10'b1111100011;
    16'b0001010010000000: out_v[150] = 10'b1010001011;
    default: out_v[150] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000000000001: out_v[151] = 10'b0010010001;
    16'b0001000000100001: out_v[151] = 10'b0101111101;
    16'b0001000000010001: out_v[151] = 10'b1011001010;
    16'b0000000000001001: out_v[151] = 10'b1011100001;
    16'b0001000000000001: out_v[151] = 10'b0000100110;
    16'b0001000000000000: out_v[151] = 10'b1001110001;
    16'b0000000000000000: out_v[151] = 10'b0001111000;
    16'b0000000000001000: out_v[151] = 10'b1011001001;
    16'b0001000000001001: out_v[151] = 10'b0100001011;
    16'b0001000000110001: out_v[151] = 10'b1001000111;
    16'b0001000000010000: out_v[151] = 10'b0001001111;
    16'b0001000000110000: out_v[151] = 10'b1000000111;
    16'b0000000000001101: out_v[151] = 10'b0101110000;
    16'b0001000000111001: out_v[151] = 10'b0100011111;
    16'b0000000000100001: out_v[151] = 10'b0010010101;
    16'b0001000000011001: out_v[151] = 10'b1000000101;
    16'b0000000000001100: out_v[151] = 10'b1101010100;
    16'b0000000000000100: out_v[151] = 10'b1011100110;
    16'b0000000000101100: out_v[151] = 10'b0110011111;
    16'b0000000000011100: out_v[151] = 10'b0000111110;
    16'b0000000000101101: out_v[151] = 10'b0001111000;
    16'b0001000000011101: out_v[151] = 10'b0101011011;
    16'b0000000000011101: out_v[151] = 10'b1111111011;
    16'b1000000000001100: out_v[151] = 10'b1111010111;
    16'b0001000000000100: out_v[151] = 10'b1001101010;
    16'b0000000000000101: out_v[151] = 10'b0100100110;
    16'b0001000000001100: out_v[151] = 10'b0011001100;
    16'b0001000000011100: out_v[151] = 10'b0101100111;
    16'b0001000000001101: out_v[151] = 10'b1101001000;
    16'b0001000000000101: out_v[151] = 10'b0010011110;
    16'b0001010000000101: out_v[151] = 10'b0010011111;
    16'b1001000000001100: out_v[151] = 10'b0111100111;
    16'b0001000000001000: out_v[151] = 10'b0111110000;
    16'b0001000000010101: out_v[151] = 10'b0100100101;
    16'b0001000000010100: out_v[151] = 10'b1010100100;
    16'b1000000000001000: out_v[151] = 10'b1000000111;
    16'b0001000000011000: out_v[151] = 10'b0000110111;
    16'b0000000000010001: out_v[151] = 10'b0111110110;
    16'b0000000000111000: out_v[151] = 10'b0100111110;
    16'b0000000000011000: out_v[151] = 10'b0000111110;
    16'b0000000000100000: out_v[151] = 10'b0000011110;
    16'b0000000000011001: out_v[151] = 10'b1010100110;
    16'b0000000000111101: out_v[151] = 10'b0000011010;
    16'b0000000000111100: out_v[151] = 10'b0111001101;
    16'b0000000000100100: out_v[151] = 10'b0100110100;
    16'b0000000000101000: out_v[151] = 10'b0010110101;
    16'b0001000000111000: out_v[151] = 10'b1111011100;
    16'b0001000000111101: out_v[151] = 10'b1101001100;
    16'b0000000000111001: out_v[151] = 10'b0000101100;
    16'b0000000000010000: out_v[151] = 10'b1110101110;
    16'b0001000000111100: out_v[151] = 10'b1110010111;
    16'b0000000000100101: out_v[151] = 10'b1000000011;
    16'b0000000000110100: out_v[151] = 10'b1011100111;
    16'b0001000000110100: out_v[151] = 10'b0110000011;
    16'b0000000000010100: out_v[151] = 10'b0110111100;
    16'b0000000000110000: out_v[151] = 10'b1111010001;
    16'b0000000000101001: out_v[151] = 10'b1011100010;
    16'b0001000000110101: out_v[151] = 10'b0101100001;
    16'b0000000000110101: out_v[151] = 10'b1101001001;
    default: out_v[151] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001000001000000: out_v[152] = 10'b0100011110;
    16'b0001101000000000: out_v[152] = 10'b1110001110;
    16'b0001101000100000: out_v[152] = 10'b1011011001;
    16'b0001111000000000: out_v[152] = 10'b0001011000;
    16'b0001000000000000: out_v[152] = 10'b0010000011;
    16'b0011100000000000: out_v[152] = 10'b1101000111;
    16'b0000101000100000: out_v[152] = 10'b0100110001;
    16'b0010101100000000: out_v[152] = 10'b0011001001;
    16'b0001101100000000: out_v[152] = 10'b1001101001;
    16'b0000101000000000: out_v[152] = 10'b1010001011;
    16'b0001001000000000: out_v[152] = 10'b1110011100;
    16'b0011101101001000: out_v[152] = 10'b0001100010;
    16'b0001001000100000: out_v[152] = 10'b0000010011;
    16'b0011000000000000: out_v[152] = 10'b0011010001;
    16'b0011101000000000: out_v[152] = 10'b0011110010;
    16'b0001101100100000: out_v[152] = 10'b0110100011;
    16'b0001100001000000: out_v[152] = 10'b1110010111;
    16'b0000101100100000: out_v[152] = 10'b1100111011;
    16'b0000001000000000: out_v[152] = 10'b1110011001;
    16'b0011101101000000: out_v[152] = 10'b0101011000;
    16'b0010111000000000: out_v[152] = 10'b0001110011;
    16'b0011100101000000: out_v[152] = 10'b0111111011;
    16'b0001111001000000: out_v[152] = 10'b1111110111;
    16'b0001100100000000: out_v[152] = 10'b0000111101;
    16'b0000011000000000: out_v[152] = 10'b1001001111;
    16'b0000001000100000: out_v[152] = 10'b0011001111;
    16'b0001100000000000: out_v[152] = 10'b1101010110;
    16'b0011101001000000: out_v[152] = 10'b0011010101;
    16'b0011101100100000: out_v[152] = 10'b0010110011;
    16'b0000101100000000: out_v[152] = 10'b0011011110;
    16'b0000111000000000: out_v[152] = 10'b1111011011;
    16'b0011101100000000: out_v[152] = 10'b1100111010;
    16'b0010111100000000: out_v[152] = 10'b1110000011;
    16'b0011111100000000: out_v[152] = 10'b0000110011;
    16'b0000000000000000: out_v[152] = 10'b1011101010;
    16'b0011100001000000: out_v[152] = 10'b0101010011;
    16'b0011111101000000: out_v[152] = 10'b0101011000;
    16'b0010101000000000: out_v[152] = 10'b0111011000;
    16'b0011100100000000: out_v[152] = 10'b1101101000;
    16'b0011111000000000: out_v[152] = 10'b1011010111;
    16'b0011111001000000: out_v[152] = 10'b0011011111;
    16'b0011100001001000: out_v[152] = 10'b0101010101;
    16'b0011100101001000: out_v[152] = 10'b1000101111;
    16'b0011111101001000: out_v[152] = 10'b0000011101;
    16'b0000100100001000: out_v[152] = 10'b0011000111;
    16'b0000100000001000: out_v[152] = 10'b0100011010;
    16'b0000100001001000: out_v[152] = 10'b0100111001;
    16'b0000000100001000: out_v[152] = 10'b0001010101;
    16'b0000000000001000: out_v[152] = 10'b0100111110;
    16'b0000100101001000: out_v[152] = 10'b0010011110;
    16'b0010100101001000: out_v[152] = 10'b1101001011;
    16'b0000100000000000: out_v[152] = 10'b0110110010;
    16'b0000000101001000: out_v[152] = 10'b1010111001;
    16'b0010100001001000: out_v[152] = 10'b1000111001;
    16'b0000010000001000: out_v[152] = 10'b1010011011;
    16'b0010100100001000: out_v[152] = 10'b1110100011;
    16'b0000000001001000: out_v[152] = 10'b0100110010;
    16'b0000100100000000: out_v[152] = 10'b0110111101;
    16'b0010100100000000: out_v[152] = 10'b0111000100;
    16'b0010101101001000: out_v[152] = 10'b1110100110;
    16'b0010100000000000: out_v[152] = 10'b0011001100;
    16'b0000110100001000: out_v[152] = 10'b1001110110;
    16'b0011100000001000: out_v[152] = 10'b1111001101;
    16'b0000100100101000: out_v[152] = 10'b0100110111;
    16'b0011101100001000: out_v[152] = 10'b0000101000;
    16'b0001100100001000: out_v[152] = 10'b0110011001;
    16'b0011111100000001: out_v[152] = 10'b0001111100;
    16'b0010110100000000: out_v[152] = 10'b0001110100;
    16'b0010101100001000: out_v[152] = 10'b1111101010;
    16'b0011001100001000: out_v[152] = 10'b1111100111;
    16'b0011100100001000: out_v[152] = 10'b0011101010;
    16'b0011101000001000: out_v[152] = 10'b1010001001;
    16'b0001100001001000: out_v[152] = 10'b0110000110;
    16'b0001100101001000: out_v[152] = 10'b0001011111;
    16'b0011001000001000: out_v[152] = 10'b1000010101;
    16'b0011001100000000: out_v[152] = 10'b1101100010;
    16'b0010100100100000: out_v[152] = 10'b0001000100;
    16'b0001101101001000: out_v[152] = 10'b1111001110;
    16'b0001101100001000: out_v[152] = 10'b0001011000;
    16'b0010100000001000: out_v[152] = 10'b1100110000;
    16'b0010100100101000: out_v[152] = 10'b0110100100;
    16'b0011110100000000: out_v[152] = 10'b1111111010;
    16'b0011001001001000: out_v[152] = 10'b0001100110;
    16'b0011111100001000: out_v[152] = 10'b1111010001;
    16'b0010000001001000: out_v[152] = 10'b0000111101;
    16'b0010110001001000: out_v[152] = 10'b0111011010;
    16'b0010110000000000: out_v[152] = 10'b1111010010;
    16'b0000110001001000: out_v[152] = 10'b1001011111;
    16'b0000110001001001: out_v[152] = 10'b0010111110;
    16'b0010000000101000: out_v[152] = 10'b1001011000;
    16'b0010110001001001: out_v[152] = 10'b1110110000;
    16'b0000000001000000: out_v[152] = 10'b1001001010;
    16'b0010000001101000: out_v[152] = 10'b1000111111;
    16'b0000100001000000: out_v[152] = 10'b0001001111;
    16'b0010110101001000: out_v[152] = 10'b0000111010;
    16'b0010100001000000: out_v[152] = 10'b0011110000;
    16'b0010010001001000: out_v[152] = 10'b1000001001;
    16'b0000010001001001: out_v[152] = 10'b1001111110;
    16'b0010000000001000: out_v[152] = 10'b1000111000;
    16'b0010010001001001: out_v[152] = 10'b0101001010;
    16'b0010000001000000: out_v[152] = 10'b0000010111;
    16'b0000000001101000: out_v[152] = 10'b0001001011;
    16'b0000010001001000: out_v[152] = 10'b1001110111;
    16'b0010000000000000: out_v[152] = 10'b1011100111;
    16'b0010110101001001: out_v[152] = 10'b0010011010;
    16'b0011000001001000: out_v[152] = 10'b0110000110;
    16'b0011001000100000: out_v[152] = 10'b1101011010;
    16'b0010000001101100: out_v[152] = 10'b0001110001;
    16'b0011000000100000: out_v[152] = 10'b1010011001;
    16'b0010000000101100: out_v[152] = 10'b1111100111;
    16'b0010000000100000: out_v[152] = 10'b0011110001;
    16'b0011001000000000: out_v[152] = 10'b0010010000;
    16'b0010000000000100: out_v[152] = 10'b1011100111;
    16'b0011000000001000: out_v[152] = 10'b1001110111;
    16'b0011001000101000: out_v[152] = 10'b0100110011;
    16'b0011101001001000: out_v[152] = 10'b0101010000;
    16'b0010000001001100: out_v[152] = 10'b1001001111;
    16'b0010000000001100: out_v[152] = 10'b1011110101;
    16'b0000100101000000: out_v[152] = 10'b0011111000;
    16'b0010101001001000: out_v[152] = 10'b1110101100;
    16'b0000000001100000: out_v[152] = 10'b1011110000;
    16'b0000101101001000: out_v[152] = 10'b1010101010;
    16'b0010100101000000: out_v[152] = 10'b1010001000;
    16'b0001100000001000: out_v[152] = 10'b1011000000;
    16'b0001101100101000: out_v[152] = 10'b0011011010;
    16'b0011100100100000: out_v[152] = 10'b1111011010;
    16'b0001100100101000: out_v[152] = 10'b1001001011;
    16'b0000000000100000: out_v[152] = 10'b0010100110;
    16'b0010100000100000: out_v[152] = 10'b0010010000;
    16'b0000100000100000: out_v[152] = 10'b1011110100;
    16'b0010000000100100: out_v[152] = 10'b0110110110;
    16'b0010100101101000: out_v[152] = 10'b1100001011;
    16'b0010000101001000: out_v[152] = 10'b0111010011;
    16'b0010100101101100: out_v[152] = 10'b0101010111;
    16'b0010000100001000: out_v[152] = 10'b0110010010;
    16'b0001000001001000: out_v[152] = 10'b0111000001;
    16'b0010000101101000: out_v[152] = 10'b0111110001;
    16'b0011000000100100: out_v[152] = 10'b1111000110;
    16'b0010100001101000: out_v[152] = 10'b1000011011;
    16'b0011000100000000: out_v[152] = 10'b1100001010;
    default: out_v[152] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0110000000100000: out_v[153] = 10'b1010100110;
    16'b0000100000111100: out_v[153] = 10'b0111110110;
    16'b1110100000111100: out_v[153] = 10'b1001001101;
    16'b0010100000111000: out_v[153] = 10'b0011111111;
    16'b0110100000100000: out_v[153] = 10'b0001010111;
    16'b0100000010110000: out_v[153] = 10'b1000111111;
    16'b0110100000101000: out_v[153] = 10'b0001101011;
    16'b0100100010001100: out_v[153] = 10'b0011011011;
    16'b0100100000001000: out_v[153] = 10'b1000011011;
    16'b0110100000111100: out_v[153] = 10'b0010110001;
    16'b0100100000101100: out_v[153] = 10'b0111110110;
    16'b0110000000110000: out_v[153] = 10'b1101001111;
    16'b0110000000111000: out_v[153] = 10'b1010101011;
    16'b0110100000110000: out_v[153] = 10'b1100001001;
    16'b0100100000001100: out_v[153] = 10'b1001101100;
    16'b0100100010011000: out_v[153] = 10'b1001001011;
    16'b0110100000111000: out_v[153] = 10'b1011101010;
    16'b0110100010110000: out_v[153] = 10'b1001111001;
    16'b0100100000111100: out_v[153] = 10'b1010011100;
    16'b0100100000110000: out_v[153] = 10'b1101101010;
    16'b0010100000101100: out_v[153] = 10'b0100001110;
    16'b0010100000001000: out_v[153] = 10'b1011010111;
    16'b0010100000111100: out_v[153] = 10'b0101110111;
    16'b0100100010111100: out_v[153] = 10'b1010110100;
    16'b0000100000110000: out_v[153] = 10'b0101001111;
    16'b0110100000010000: out_v[153] = 10'b1111101110;
    16'b0000100000101100: out_v[153] = 10'b0101111011;
    16'b0010100000101000: out_v[153] = 10'b0001000001;
    16'b0110100000101100: out_v[153] = 10'b1110111110;
    16'b0100100010111000: out_v[153] = 10'b0110010011;
    16'b0100100010011100: out_v[153] = 10'b1010111110;
    16'b0110000010110000: out_v[153] = 10'b0111000101;
    16'b0000100000111000: out_v[153] = 10'b1101111010;
    16'b0010100000110000: out_v[153] = 10'b1110110111;
    16'b0100010010100000: out_v[153] = 10'b1100101001;
    16'b0100100010110000: out_v[153] = 10'b1000111011;
    16'b0100000010100000: out_v[153] = 10'b0100011011;
    16'b0000100000110100: out_v[153] = 10'b0011011101;
    16'b0110100010111000: out_v[153] = 10'b1100100111;
    16'b0110100010111100: out_v[153] = 10'b0111011000;
    16'b0100110010011100: out_v[153] = 10'b1010111011;
    16'b0100100000111000: out_v[153] = 10'b0011111111;
    16'b0100010000000000: out_v[153] = 10'b0011001010;
    16'b0100000000000000: out_v[153] = 10'b0111100110;
    16'b0000000000000000: out_v[153] = 10'b1010110010;
    16'b0000010000100000: out_v[153] = 10'b1100111011;
    16'b0000000000100000: out_v[153] = 10'b0101101010;
    16'b0000010000000000: out_v[153] = 10'b1001011101;
    16'b0010000000100000: out_v[153] = 10'b0101100110;
    16'b0010010000100000: out_v[153] = 10'b0001001010;
    16'b0000000010100000: out_v[153] = 10'b1110011000;
    16'b0110000010100000: out_v[153] = 10'b1101010110;
    16'b0100000010010000: out_v[153] = 10'b1010011011;
    16'b0100010010001000: out_v[153] = 10'b0100000110;
    16'b0100000010011000: out_v[153] = 10'b0111001111;
    16'b0100110010001100: out_v[153] = 10'b0011001110;
    16'b0000000010000000: out_v[153] = 10'b0111000110;
    16'b0110010000110000: out_v[153] = 10'b0011010100;
    16'b0110100010100000: out_v[153] = 10'b0101010110;
    16'b0100010010000000: out_v[153] = 10'b0010101101;
    16'b0110000010011000: out_v[153] = 10'b1111011011;
    16'b0110100010011000: out_v[153] = 10'b0101111000;
    16'b0100000000100000: out_v[153] = 10'b1110000101;
    16'b0000010010011000: out_v[153] = 10'b1101100111;
    16'b0110000000100010: out_v[153] = 10'b1111011000;
    16'b0100010010011000: out_v[153] = 10'b1111000111;
    16'b0110010000100000: out_v[153] = 10'b0010110111;
    16'b0100110010011000: out_v[153] = 10'b1111110110;
    16'b0110000010111000: out_v[153] = 10'b1001110000;
    16'b0100000010000000: out_v[153] = 10'b1001101010;
    16'b0110000000000000: out_v[153] = 10'b1000110101;
    16'b0100110010001000: out_v[153] = 10'b0000100110;
    16'b0110000010000000: out_v[153] = 10'b1101011110;
    16'b0100000010001000: out_v[153] = 10'b0111011100;
    16'b0000000010011000: out_v[153] = 10'b0110011010;
    16'b0000000010010000: out_v[153] = 10'b0110010111;
    16'b0000010010010000: out_v[153] = 10'b0100010100;
    16'b0010000010100000: out_v[153] = 10'b1001001110;
    16'b0100000000010000: out_v[153] = 10'b1001010101;
    16'b0100010000010000: out_v[153] = 10'b0011000110;
    16'b0100010010010000: out_v[153] = 10'b0101000111;
    16'b0110010000111000: out_v[153] = 10'b1001001111;
    16'b0110100010011100: out_v[153] = 10'b1011111010;
    16'b0010010010100000: out_v[153] = 10'b0001010011;
    16'b0000010010100000: out_v[153] = 10'b0000011101;
    16'b0010010010000000: out_v[153] = 10'b0010011001;
    16'b0010000010000000: out_v[153] = 10'b1101011011;
    16'b0010010000000000: out_v[153] = 10'b1100001010;
    16'b0010011000100000: out_v[153] = 10'b1101000111;
    16'b0010110010100100: out_v[153] = 10'b0011101011;
    16'b0010011010100000: out_v[153] = 10'b1000001010;
    16'b0100010000100000: out_v[153] = 10'b0111011000;
    16'b0000010010000000: out_v[153] = 10'b1001011101;
    16'b0010000000000000: out_v[153] = 10'b0110101000;
    16'b0110010010100000: out_v[153] = 10'b1000111000;
    16'b0010001000100000: out_v[153] = 10'b1110010110;
    16'b0000110010100000: out_v[153] = 10'b1001011011;
    16'b0110000000101000: out_v[153] = 10'b1110111110;
    16'b0000110010100100: out_v[153] = 10'b0101011111;
    16'b0010110010100000: out_v[153] = 10'b1000101111;
    16'b0100110010000100: out_v[153] = 10'b1001011001;
    16'b0110011010100000: out_v[153] = 10'b1011111001;
    16'b0000000010001000: out_v[153] = 10'b0001010110;
    16'b0010000010111000: out_v[153] = 10'b0010011000;
    16'b0000110010000100: out_v[153] = 10'b1011011101;
    16'b0010000010011000: out_v[153] = 10'b0111011010;
    16'b0000100010000100: out_v[153] = 10'b1101011100;
    16'b0010100010111100: out_v[153] = 10'b1010110110;
    16'b0010000010010000: out_v[153] = 10'b0110011000;
    16'b0000000010111000: out_v[153] = 10'b1001011010;
    16'b0010010010111000: out_v[153] = 10'b1000111000;
    16'b0010000010110000: out_v[153] = 10'b1011100100;
    16'b0000000010110000: out_v[153] = 10'b1000011010;
    16'b0000100010111100: out_v[153] = 10'b0100011111;
    16'b0000100010011100: out_v[153] = 10'b1000000111;
    16'b0010000000100100: out_v[153] = 10'b1110110111;
    16'b0000010010100100: out_v[153] = 10'b0011110111;
    16'b1100110000000100: out_v[153] = 10'b0000110111;
    16'b1100010000000100: out_v[153] = 10'b1010110111;
    16'b0010010010100100: out_v[153] = 10'b1101010011;
    16'b1010010010100100: out_v[153] = 10'b1101111010;
    16'b0100000000111000: out_v[153] = 10'b1010011100;
    16'b0110010010110000: out_v[153] = 10'b1101110010;
    16'b0100010010110000: out_v[153] = 10'b0001010110;
    16'b0010000000110000: out_v[153] = 10'b0011101011;
    16'b0100010000110000: out_v[153] = 10'b1110110100;
    16'b0110110000110000: out_v[153] = 10'b0011010101;
    16'b0100000010111000: out_v[153] = 10'b0010111100;
    16'b0110010010111000: out_v[153] = 10'b1001011011;
    16'b0100000000011000: out_v[153] = 10'b0111101000;
    16'b0100000000110000: out_v[153] = 10'b1011010100;
    16'b1000100010000100: out_v[153] = 10'b0011011011;
    16'b0010100000100000: out_v[153] = 10'b1001100010;
    16'b0000100010000000: out_v[153] = 10'b1110000010;
    16'b0000100010100100: out_v[153] = 10'b1011011000;
    16'b0000100000000100: out_v[153] = 10'b0011100111;
    16'b0000100010100000: out_v[153] = 10'b1010100101;
    16'b0100100000000100: out_v[153] = 10'b0011100110;
    16'b0010100010100000: out_v[153] = 10'b0011101000;
    16'b1100100010000100: out_v[153] = 10'b0111011010;
    16'b0100100010000000: out_v[153] = 10'b0110010010;
    16'b0100100010000100: out_v[153] = 10'b0110110010;
    16'b0100100000000000: out_v[153] = 10'b0000100010;
    16'b0000100000000000: out_v[153] = 10'b1000101001;
    16'b0100110000100000: out_v[153] = 10'b0111000010;
    16'b0110110000100000: out_v[153] = 10'b1000011000;
    16'b0110110010100100: out_v[153] = 10'b0100111000;
    16'b0100110000000100: out_v[153] = 10'b1100101000;
    16'b0100110000100100: out_v[153] = 10'b1010001101;
    16'b0000110000100100: out_v[153] = 10'b0011011011;
    16'b1110110010100100: out_v[153] = 10'b0001101110;
    16'b1000110000000100: out_v[153] = 10'b1101000111;
    16'b1000110000010100: out_v[153] = 10'b0111001111;
    16'b0110010010000000: out_v[153] = 10'b0110000000;
    16'b0000110000000100: out_v[153] = 10'b1001101010;
    16'b0100110000000000: out_v[153] = 10'b1100101010;
    16'b0100110010100000: out_v[153] = 10'b0111110001;
    16'b0000110000010100: out_v[153] = 10'b1110101011;
    16'b0100100000100000: out_v[153] = 10'b0110011010;
    16'b0110110000100100: out_v[153] = 10'b1011111110;
    16'b1100110000100100: out_v[153] = 10'b1011010111;
    16'b0100110010100100: out_v[153] = 10'b0010001100;
    16'b0110010000000000: out_v[153] = 10'b1110101011;
    16'b0110110010100000: out_v[153] = 10'b0100111001;
    16'b0000100010111000: out_v[153] = 10'b0010111111;
    16'b0000110000000000: out_v[153] = 10'b1011001011;
    16'b0000110010000000: out_v[153] = 10'b1000010111;
    16'b0010100010111000: out_v[153] = 10'b0011001010;
    16'b0000100010010000: out_v[153] = 10'b1101111011;
    default: out_v[153] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1010000100001000: out_v[154] = 10'b1010111011;
    16'b1010000000001000: out_v[154] = 10'b1000100011;
    16'b0010000000001000: out_v[154] = 10'b1101100011;
    16'b0001000100000000: out_v[154] = 10'b1011101011;
    16'b0001000000001000: out_v[154] = 10'b1010001110;
    16'b1001000000001000: out_v[154] = 10'b0111011101;
    16'b1001000100001000: out_v[154] = 10'b1001011011;
    16'b1010000000011000: out_v[154] = 10'b0101101011;
    16'b0001000000000000: out_v[154] = 10'b1000110111;
    16'b1000000000001000: out_v[154] = 10'b1011000001;
    16'b1010000000101000: out_v[154] = 10'b1011001110;
    16'b1000000100001000: out_v[154] = 10'b1111001000;
    16'b0010000100001000: out_v[154] = 10'b0100011000;
    16'b0000000000001000: out_v[154] = 10'b1000101110;
    16'b1011000100001000: out_v[154] = 10'b0011111010;
    16'b1011001100001000: out_v[154] = 10'b0110110001;
    16'b1011001100000000: out_v[154] = 10'b0010110011;
    16'b0001001100000000: out_v[154] = 10'b0010011001;
    16'b1001000100000000: out_v[154] = 10'b0100100111;
    16'b0000000000011000: out_v[154] = 10'b1000010111;
    16'b1000000000000000: out_v[154] = 10'b0110101000;
    16'b1001001100001000: out_v[154] = 10'b0011011111;
    16'b1001000100011000: out_v[154] = 10'b1011101110;
    16'b0010000000011000: out_v[154] = 10'b0100110001;
    16'b1000000000011000: out_v[154] = 10'b0011011011;
    16'b1010000000000000: out_v[154] = 10'b0000100011;
    16'b0001000100001000: out_v[154] = 10'b0111001000;
    16'b0011000100001000: out_v[154] = 10'b0001001001;
    16'b1001001100000000: out_v[154] = 10'b1110010011;
    16'b0010000000000000: out_v[154] = 10'b1110011011;
    16'b1010000100000000: out_v[154] = 10'b1100100110;
    16'b1001000000011000: out_v[154] = 10'b1100111111;
    16'b1000000100000000: out_v[154] = 10'b1100010101;
    16'b1011000100000000: out_v[154] = 10'b0100110010;
    16'b0000000000100000: out_v[154] = 10'b1011100001;
    16'b1000000000100000: out_v[154] = 10'b0110101111;
    16'b0000000000000000: out_v[154] = 10'b1111100110;
    16'b0000000100100000: out_v[154] = 10'b0101001111;
    16'b0000000000110000: out_v[154] = 10'b0111011001;
    16'b1000000100100000: out_v[154] = 10'b1010110111;
    16'b1011000000101000: out_v[154] = 10'b1010110100;
    16'b1001000100100000: out_v[154] = 10'b0011101010;
    16'b1001000100110000: out_v[154] = 10'b1111101100;
    16'b1010000000100000: out_v[154] = 10'b0111001010;
    16'b1011000000100000: out_v[154] = 10'b1000101101;
    16'b0001000000100000: out_v[154] = 10'b0010100010;
    16'b1010000100010000: out_v[154] = 10'b1100100100;
    16'b1010000100100000: out_v[154] = 10'b0111001011;
    16'b1010000000010000: out_v[154] = 10'b1111001010;
    16'b1010000100110000: out_v[154] = 10'b0001111001;
    16'b1001000000100000: out_v[154] = 10'b1000000110;
    16'b1010000100101000: out_v[154] = 10'b1101100110;
    16'b1001000000101000: out_v[154] = 10'b0011010100;
    16'b1000000100110000: out_v[154] = 10'b0001010111;
    16'b0011000000100000: out_v[154] = 10'b0101110111;
    16'b1001000000000000: out_v[154] = 10'b1000000100;
    16'b1011000100100000: out_v[154] = 10'b1001111011;
    16'b1011000000000000: out_v[154] = 10'b0110001100;
    16'b0010000100100000: out_v[154] = 10'b1001001010;
    16'b1001000000110000: out_v[154] = 10'b1011110100;
    16'b0010000000100000: out_v[154] = 10'b0111010001;
    16'b1011000000110000: out_v[154] = 10'b0100111110;
    16'b1010000000110000: out_v[154] = 10'b0101100000;
    16'b0001000100100000: out_v[154] = 10'b1001100110;
    16'b0010000000110000: out_v[154] = 10'b0111001010;
    16'b1011000100110000: out_v[154] = 10'b0011001011;
    16'b1000000100101000: out_v[154] = 10'b0000001110;
    16'b1000000000110000: out_v[154] = 10'b0000010011;
    16'b1000000000101000: out_v[154] = 10'b0000111000;
    16'b0000000100101000: out_v[154] = 10'b0001110011;
    16'b0000000001100000: out_v[154] = 10'b1101101100;
    16'b0010000100000000: out_v[154] = 10'b1000011110;
    16'b1000000000111000: out_v[154] = 10'b0010110011;
    16'b1010000100011000: out_v[154] = 10'b1100011011;
    16'b1001000100101000: out_v[154] = 10'b0011111011;
    16'b1011000100011000: out_v[154] = 10'b1011101000;
    16'b1000000000010000: out_v[154] = 10'b0111010111;
    16'b1010000000111000: out_v[154] = 10'b1000100111;
    16'b0011000100000000: out_v[154] = 10'b0101111010;
    16'b0001000100101000: out_v[154] = 10'b1001101011;
    16'b0000000100000000: out_v[154] = 10'b1000100101;
    16'b1011000100101000: out_v[154] = 10'b1111000111;
    16'b0000000101100000: out_v[154] = 10'b0110011010;
    16'b1011000100010000: out_v[154] = 10'b0111001010;
    16'b1000000100111000: out_v[154] = 10'b0011100111;
    16'b0010000000101000: out_v[154] = 10'b0001011100;
    16'b0010000001101000: out_v[154] = 10'b0110000110;
    16'b0000000000101000: out_v[154] = 10'b1000110010;
    16'b0010000100101000: out_v[154] = 10'b0000011101;
    16'b0010001100101000: out_v[154] = 10'b0101010111;
    16'b0010001000101000: out_v[154] = 10'b0110001110;
    16'b0000000001101000: out_v[154] = 10'b1001101011;
    16'b0010001100100000: out_v[154] = 10'b1000011110;
    16'b0001000000101000: out_v[154] = 10'b0000111111;
    16'b0010001000100000: out_v[154] = 10'b1011111001;
    16'b0000000000111000: out_v[154] = 10'b0111100011;
    16'b0000000001001000: out_v[154] = 10'b1000100110;
    16'b0000000100001000: out_v[154] = 10'b0111100010;
    16'b0000000101101000: out_v[154] = 10'b0010101110;
    16'b0011000100101000: out_v[154] = 10'b1001110110;
    16'b0011000000101000: out_v[154] = 10'b0101110110;
    16'b0011000000001000: out_v[154] = 10'b1011001010;
    16'b0010000001001000: out_v[154] = 10'b0110000110;
    16'b0010001100000000: out_v[154] = 10'b1111111010;
    16'b0010000001000000: out_v[154] = 10'b0111110110;
    16'b0010000001100000: out_v[154] = 10'b0101000100;
    16'b0010001000000000: out_v[154] = 10'b1100110110;
    16'b0010001001000000: out_v[154] = 10'b0111110011;
    16'b0010001001101000: out_v[154] = 10'b1011001011;
    16'b0010001100001000: out_v[154] = 10'b0110010111;
    16'b0010001001001000: out_v[154] = 10'b1000001111;
    16'b0010001001100000: out_v[154] = 10'b1100110000;
    16'b0000000001000000: out_v[154] = 10'b0001111010;
    16'b0000001000100000: out_v[154] = 10'b1011000110;
    16'b0010001000001000: out_v[154] = 10'b1110000100;
    default: out_v[154] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000001011000: out_v[155] = 10'b1000101100;
    16'b0000000010000000: out_v[155] = 10'b0100001010;
    16'b0000000001001010: out_v[155] = 10'b1100101000;
    16'b0000010001001010: out_v[155] = 10'b0001101001;
    16'b0000000001001000: out_v[155] = 10'b0001101011;
    16'b0000000010010000: out_v[155] = 10'b1000001001;
    16'b0000000011001010: out_v[155] = 10'b1001001101;
    16'b0000000000000000: out_v[155] = 10'b0001111110;
    16'b0000000000000010: out_v[155] = 10'b0100110101;
    16'b0000000001100000: out_v[155] = 10'b0000110111;
    16'b0000000011010000: out_v[155] = 10'b0011010010;
    16'b0000000000001000: out_v[155] = 10'b0001101011;
    16'b0000010000001000: out_v[155] = 10'b1010100010;
    16'b0000000001101010: out_v[155] = 10'b0100111011;
    16'b0000000011001000: out_v[155] = 10'b0110111101;
    16'b0000000001000000: out_v[155] = 10'b0001111011;
    16'b0000000001010000: out_v[155] = 10'b0110001001;
    16'b0000000011011010: out_v[155] = 10'b1110100010;
    16'b0000000011101010: out_v[155] = 10'b0100001011;
    16'b0000000000010000: out_v[155] = 10'b1111010010;
    16'b0000000011011000: out_v[155] = 10'b1011001011;
    16'b0000000001101000: out_v[155] = 10'b1000100101;
    16'b0000000010001000: out_v[155] = 10'b1011100100;
    16'b0000000001100010: out_v[155] = 10'b1110010011;
    16'b0000000001000010: out_v[155] = 10'b1101101001;
    16'b0000000001011010: out_v[155] = 10'b1001000010;
    16'b0000010000000000: out_v[155] = 10'b0111100111;
    16'b0000010000010000: out_v[155] = 10'b1011110111;
    16'b0000000011101000: out_v[155] = 10'b0010001011;
    16'b0000010010010000: out_v[155] = 10'b0011011010;
    16'b0000000000001010: out_v[155] = 10'b0111010110;
    16'b0000000011111000: out_v[155] = 10'b0101110101;
    16'b0000000000011000: out_v[155] = 10'b1011001001;
    16'b0000000011111010: out_v[155] = 10'b1010000101;
    16'b0000010011001010: out_v[155] = 10'b1010011100;
    16'b0000000011000010: out_v[155] = 10'b1010110110;
    16'b0000000011100010: out_v[155] = 10'b1010100111;
    16'b0000000011000000: out_v[155] = 10'b0001010100;
    16'b0000000011100000: out_v[155] = 10'b0101010000;
    16'b0000000010101000: out_v[155] = 10'b0010101000;
    16'b0000000001110000: out_v[155] = 10'b0011111000;
    16'b0000000010110000: out_v[155] = 10'b1101000110;
    16'b0000000011110000: out_v[155] = 10'b0010000110;
    16'b0000000010111000: out_v[155] = 10'b0010011001;
    16'b0000000010100000: out_v[155] = 10'b0011001100;
    16'b0000010001011000: out_v[155] = 10'b0011111101;
    16'b0000000000110000: out_v[155] = 10'b1110001110;
    16'b0000010010001000: out_v[155] = 10'b1000000101;
    16'b0000000010011000: out_v[155] = 10'b1001110001;
    16'b0000000000101000: out_v[155] = 10'b1111000111;
    16'b0000010000010100: out_v[155] = 10'b0110001111;
    16'b0000000001111000: out_v[155] = 10'b0100100111;
    16'b0000000000100000: out_v[155] = 10'b1101001101;
    16'b0000010001111000: out_v[155] = 10'b0011011111;
    16'b0000010001010000: out_v[155] = 10'b0000111110;
    16'b0000000000111000: out_v[155] = 10'b1101000101;
    16'b0000010000011000: out_v[155] = 10'b1011011010;
    16'b0000010011001000: out_v[155] = 10'b1100100100;
    16'b0000010010010100: out_v[155] = 10'b1101011111;
    16'b0000010011010100: out_v[155] = 10'b0011001110;
    16'b0000010011010000: out_v[155] = 10'b0111011111;
    16'b0000010011111000: out_v[155] = 10'b1001001111;
    16'b0000010011111100: out_v[155] = 10'b0111110111;
    16'b0000000010010010: out_v[155] = 10'b0010011001;
    16'b0000000011010010: out_v[155] = 10'b1000000001;
    16'b0000000001010010: out_v[155] = 10'b1111110101;
    16'b0000000011110010: out_v[155] = 10'b0100010110;
    16'b0000000010011010: out_v[155] = 10'b0001110000;
    16'b0000000001111010: out_v[155] = 10'b1100110000;
    16'b0000000010000010: out_v[155] = 10'b1111100010;
    16'b0000000000010010: out_v[155] = 10'b1101010011;
    16'b0000000000011010: out_v[155] = 10'b0101011000;
    16'b0000000001110010: out_v[155] = 10'b0101100000;
    16'b0000000001011001: out_v[155] = 10'b0100110011;
    16'b0000000001111001: out_v[155] = 10'b0011110000;
    16'b0000000010101010: out_v[155] = 10'b1111001010;
    16'b0000000011101001: out_v[155] = 10'b0100011111;
    16'b0000000011001001: out_v[155] = 10'b1010111111;
    16'b0000000010001010: out_v[155] = 10'b0011011011;
    16'b0000001010010000: out_v[155] = 10'b1011001011;
    default: out_v[155] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1000001100010000: out_v[156] = 10'b1001010101;
    16'b1010001100010101: out_v[156] = 10'b0011101111;
    16'b1010000100000101: out_v[156] = 10'b0011001111;
    16'b1010001000000101: out_v[156] = 10'b1011110100;
    16'b0010001100010000: out_v[156] = 10'b0111111011;
    16'b1110000000000101: out_v[156] = 10'b0000001101;
    16'b1010001100010100: out_v[156] = 10'b1000001111;
    16'b0110000100000101: out_v[156] = 10'b1101010110;
    16'b1010000000000101: out_v[156] = 10'b1101010000;
    16'b1010001100010000: out_v[156] = 10'b1010101000;
    16'b1010001100010001: out_v[156] = 10'b0110101000;
    16'b0010000000000101: out_v[156] = 10'b0001000011;
    16'b0010000100000101: out_v[156] = 10'b1000010111;
    16'b1010001100000101: out_v[156] = 10'b1011110010;
    16'b1010000100010101: out_v[156] = 10'b1010010111;
    16'b0010000100000001: out_v[156] = 10'b1001011001;
    16'b1010001000010000: out_v[156] = 10'b0010111010;
    16'b1000001000010000: out_v[156] = 10'b1001000111;
    16'b1010001000010100: out_v[156] = 10'b1001010011;
    16'b1010000000010101: out_v[156] = 10'b1111000010;
    16'b0010000100010101: out_v[156] = 10'b1000010111;
    16'b1010001000010101: out_v[156] = 10'b0101011001;
    16'b0110000000000101: out_v[156] = 10'b1111011100;
    16'b1110000100000101: out_v[156] = 10'b1010100111;
    16'b0010001100010100: out_v[156] = 10'b0011001101;
    16'b1110001000000101: out_v[156] = 10'b1011000011;
    16'b1010001100000000: out_v[156] = 10'b0110111000;
    16'b1110000000000001: out_v[156] = 10'b1110000011;
    16'b0010001100010101: out_v[156] = 10'b0010100101;
    16'b1000001100000000: out_v[156] = 10'b0110000011;
    16'b1010000100000001: out_v[156] = 10'b1010110111;
    16'b1000000000000101: out_v[156] = 10'b1000000111;
    16'b1000000100000101: out_v[156] = 10'b1000011011;
    16'b1010000000000001: out_v[156] = 10'b0101000110;
    16'b1110001100000101: out_v[156] = 10'b1000111011;
    16'b1010001000000001: out_v[156] = 10'b0110111011;
    16'b0010001100000000: out_v[156] = 10'b0110001101;
    16'b0010000000000000: out_v[156] = 10'b0010100110;
    16'b0000000000000000: out_v[156] = 10'b0110101001;
    16'b1000000000000000: out_v[156] = 10'b0001111110;
    16'b0000000100000000: out_v[156] = 10'b1100100001;
    16'b1000000100000000: out_v[156] = 10'b0111000010;
    16'b0010000100000000: out_v[156] = 10'b0111100100;
    16'b1010000000000000: out_v[156] = 10'b0010010100;
    16'b0010001000010001: out_v[156] = 10'b1110110110;
    16'b0010001000000000: out_v[156] = 10'b0000010100;
    16'b0010001000010000: out_v[156] = 10'b1000101100;
    16'b0110000000000000: out_v[156] = 10'b0111101011;
    16'b0010001000010100: out_v[156] = 10'b1110011001;
    16'b1010000100000000: out_v[156] = 10'b1100110100;
    16'b0110000000000001: out_v[156] = 10'b1010111111;
    16'b0100000000000000: out_v[156] = 10'b1110100101;
    16'b0110001000010000: out_v[156] = 10'b1100111100;
    16'b1000001000000000: out_v[156] = 10'b1101001111;
    16'b0010000000010001: out_v[156] = 10'b1100001100;
    16'b0010001000000100: out_v[156] = 10'b0100000111;
    16'b0010001010000000: out_v[156] = 10'b0000100111;
    16'b0000001000010000: out_v[156] = 10'b1000110110;
    16'b1010001000000000: out_v[156] = 10'b0000011111;
    16'b0110001000000000: out_v[156] = 10'b1101110011;
    16'b0110001000010001: out_v[156] = 10'b1101110111;
    16'b0110000000010001: out_v[156] = 10'b1100100111;
    16'b0000001000000000: out_v[156] = 10'b1111000000;
    16'b0110000100000000: out_v[156] = 10'b1011000010;
    16'b0110000100000001: out_v[156] = 10'b0010100111;
    16'b1000001110010000: out_v[156] = 10'b0010110111;
    16'b1000000100010000: out_v[156] = 10'b0101011010;
    16'b0000000100010000: out_v[156] = 10'b0101110000;
    16'b1110001100000001: out_v[156] = 10'b1100101010;
    16'b1010000100010000: out_v[156] = 10'b0100101000;
    16'b1100001100010001: out_v[156] = 10'b1111001111;
    16'b1110001100010001: out_v[156] = 10'b1111011010;
    16'b1000001100010100: out_v[156] = 10'b0011110110;
    16'b1000001100010001: out_v[156] = 10'b0111001010;
    16'b1010001100000001: out_v[156] = 10'b1100111001;
    16'b1000000110000000: out_v[156] = 10'b1100110111;
    16'b0000001100010000: out_v[156] = 10'b0110001011;
    16'b1000000000010000: out_v[156] = 10'b0010101010;
    16'b0000001100000000: out_v[156] = 10'b0010010000;
    16'b1000001100000100: out_v[156] = 10'b0101001011;
    16'b0000000000010100: out_v[156] = 10'b0101100110;
    16'b1000001000010101: out_v[156] = 10'b1100011101;
    16'b0000000000000100: out_v[156] = 10'b1100110010;
    16'b0000001100010100: out_v[156] = 10'b1000010011;
    16'b0000001000010100: out_v[156] = 10'b1011011000;
    16'b0000001000000100: out_v[156] = 10'b1101000100;
    16'b1000001000000100: out_v[156] = 10'b0111011101;
    16'b0000000100000100: out_v[156] = 10'b1100101110;
    16'b0000001000010101: out_v[156] = 10'b0010010110;
    16'b1000001000010100: out_v[156] = 10'b0011010001;
    16'b0000001100000100: out_v[156] = 10'b0101001111;
    16'b0000000000010101: out_v[156] = 10'b1101011101;
    16'b0000000000010000: out_v[156] = 10'b0010011100;
    16'b0000001100010101: out_v[156] = 10'b0110011111;
    16'b0000000100010101: out_v[156] = 10'b0110000011;
    16'b1000000000000100: out_v[156] = 10'b0111100101;
    16'b1000001100010101: out_v[156] = 10'b0100011110;
    16'b1000000000010101: out_v[156] = 10'b1000011011;
    16'b0011000100000000: out_v[156] = 10'b1011101111;
    16'b0010000100010000: out_v[156] = 10'b1100101001;
    16'b1000000100000100: out_v[156] = 10'b0010111010;
    16'b1010000100000100: out_v[156] = 10'b0011101010;
    16'b1010000000000100: out_v[156] = 10'b1001111011;
    16'b0010000100000100: out_v[156] = 10'b1001001110;
    16'b0000001000000001: out_v[156] = 10'b1001100010;
    16'b0100001000010101: out_v[156] = 10'b1111101011;
    16'b0010001100000101: out_v[156] = 10'b0111011110;
    16'b0000001100010001: out_v[156] = 10'b0010101011;
    16'b0010001000000101: out_v[156] = 10'b0011010010;
    16'b0110001000010101: out_v[156] = 10'b1110011001;
    16'b0100001000000101: out_v[156] = 10'b0110111011;
    16'b0000001000000101: out_v[156] = 10'b0001001011;
    16'b0010001000010101: out_v[156] = 10'b0111010011;
    16'b0110001000000101: out_v[156] = 10'b0111000011;
    16'b0010001100000001: out_v[156] = 10'b0001101110;
    16'b0010001100010001: out_v[156] = 10'b1100101100;
    16'b0010001000000001: out_v[156] = 10'b1001100101;
    16'b0000001000010001: out_v[156] = 10'b1011100010;
    16'b0100001000000001: out_v[156] = 10'b1110101011;
    16'b0000001100000001: out_v[156] = 10'b0011110100;
    16'b1000011000010000: out_v[156] = 10'b0010100010;
    16'b0000011000010000: out_v[156] = 10'b1010110000;
    16'b1000011100000000: out_v[156] = 10'b1111011111;
    16'b1000011000000000: out_v[156] = 10'b1001001110;
    16'b1000010100000000: out_v[156] = 10'b1001000110;
    16'b1000010000000000: out_v[156] = 10'b0011001001;
    16'b1000011000010100: out_v[156] = 10'b1101111111;
    16'b0000010000000000: out_v[156] = 10'b0010101001;
    16'b1000011100010000: out_v[156] = 10'b0110011101;
    16'b1000011100010100: out_v[156] = 10'b0111001110;
    16'b1000000000010001: out_v[156] = 10'b1011100000;
    16'b1000001000010001: out_v[156] = 10'b0110010110;
    16'b0000011000000000: out_v[156] = 10'b1101011011;
    16'b1000011000000100: out_v[156] = 10'b1110101101;
    16'b0000001000110100: out_v[156] = 10'b1011000111;
    default: out_v[156] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100001100001000: out_v[157] = 10'b1101011011;
    16'b0100101100011010: out_v[157] = 10'b1100110010;
    16'b0100101000010010: out_v[157] = 10'b0101011000;
    16'b0100001100011010: out_v[157] = 10'b1010100011;
    16'b0100000000011010: out_v[157] = 10'b1110000001;
    16'b0000101000010010: out_v[157] = 10'b0111110111;
    16'b0000101100000010: out_v[157] = 10'b1011011100;
    16'b0100001110011000: out_v[157] = 10'b1001011001;
    16'b0100100010010000: out_v[157] = 10'b1000001111;
    16'b0100001110011010: out_v[157] = 10'b1011101010;
    16'b0100101100010010: out_v[157] = 10'b0011010101;
    16'b0100101100000010: out_v[157] = 10'b1011001111;
    16'b0100001100011000: out_v[157] = 10'b0100011010;
    16'b0000101100000000: out_v[157] = 10'b0011011001;
    16'b0000101000000000: out_v[157] = 10'b1000100111;
    16'b0000101100011010: out_v[157] = 10'b1101001111;
    16'b0000001100011010: out_v[157] = 10'b0010100110;
    16'b0100101110011000: out_v[157] = 10'b0110111111;
    16'b0100000100011010: out_v[157] = 10'b1010001111;
    16'b0100101000000010: out_v[157] = 10'b1100000001;
    16'b0100101100010000: out_v[157] = 10'b0010110101;
    16'b0000001000000000: out_v[157] = 10'b0100111000;
    16'b0000101000011010: out_v[157] = 10'b1010000110;
    16'b0100001000000010: out_v[157] = 10'b1000110101;
    16'b0100101100000000: out_v[157] = 10'b1010001111;
    16'b0100001000011010: out_v[157] = 10'b0010100110;
    16'b0000101100001000: out_v[157] = 10'b1111100010;
    16'b0000101000010000: out_v[157] = 10'b0010100011;
    16'b0000101100010010: out_v[157] = 10'b1110110110;
    16'b0100101110011010: out_v[157] = 10'b1111100001;
    16'b0100101000010000: out_v[157] = 10'b1000011111;
    16'b0100000110011010: out_v[157] = 10'b0011000011;
    16'b0000001000000010: out_v[157] = 10'b0111100001;
    16'b0100101010000010: out_v[157] = 10'b0111011011;
    16'b0100101000011010: out_v[157] = 10'b0111100111;
    16'b0000001100011000: out_v[157] = 10'b1000000111;
    16'b0100101100011000: out_v[157] = 10'b0101010100;
    16'b0000001100001000: out_v[157] = 10'b1101000111;
    16'b0100101000000000: out_v[157] = 10'b0100110010;
    16'b0000101000000010: out_v[157] = 10'b1110100101;
    16'b0000101100010000: out_v[157] = 10'b0000001001;
    16'b0100101010011010: out_v[157] = 10'b0101111010;
    16'b0100101010010010: out_v[157] = 10'b1011110110;
    16'b0100101110010010: out_v[157] = 10'b0010100111;
    16'b0100101110010000: out_v[157] = 10'b0101010100;
    16'b0100101100001000: out_v[157] = 10'b1101001010;
    16'b0000101100011000: out_v[157] = 10'b0001100100;
    16'b0000000010000010: out_v[157] = 10'b1000110111;
    16'b0000000010010010: out_v[157] = 10'b0001011111;
    16'b0100001010010000: out_v[157] = 10'b1001110110;
    16'b0100000000010000: out_v[157] = 10'b1101101011;
    16'b0100001000010000: out_v[157] = 10'b0110010111;
    16'b0000000010000000: out_v[157] = 10'b1000110011;
    16'b0100000010000000: out_v[157] = 10'b0011111000;
    16'b0100001010000000: out_v[157] = 10'b1110010001;
    16'b0100000010010000: out_v[157] = 10'b0001100101;
    16'b0100000010000010: out_v[157] = 10'b0000011111;
    16'b0100001000000000: out_v[157] = 10'b0100011010;
    16'b0000000010010000: out_v[157] = 10'b0001110101;
    16'b0100000000000000: out_v[157] = 10'b1111101111;
    16'b0000000110000010: out_v[157] = 10'b1011010110;
    16'b0100001010010010: out_v[157] = 10'b0101111001;
    16'b0000001010010000: out_v[157] = 10'b1110001101;
    16'b0000001010000000: out_v[157] = 10'b1001000110;
    16'b0100101010010000: out_v[157] = 10'b1000011110;
    16'b0000101110001000: out_v[157] = 10'b0100010010;
    16'b0000001110000000: out_v[157] = 10'b1110001111;
    16'b0000001000011000: out_v[157] = 10'b0111100111;
    16'b0000001010011000: out_v[157] = 10'b1000011000;
    16'b0000001000011010: out_v[157] = 10'b1110000000;
    16'b0000001110010000: out_v[157] = 10'b1110000101;
    16'b0000101110011000: out_v[157] = 10'b1111000110;
    16'b0000000100011010: out_v[157] = 10'b0110100011;
    16'b0100001010011000: out_v[157] = 10'b0010111101;
    16'b0000101100001010: out_v[157] = 10'b1011001111;
    16'b0000001100001010: out_v[157] = 10'b1111101011;
    16'b0000101010010000: out_v[157] = 10'b1101110110;
    16'b0000101000011000: out_v[157] = 10'b0011110100;
    16'b0000101110010010: out_v[157] = 10'b1001110111;
    16'b0000101110000000: out_v[157] = 10'b0001101110;
    16'b0000101010011000: out_v[157] = 10'b0010111011;
    16'b0000101010010010: out_v[157] = 10'b1001011001;
    16'b0000001100000010: out_v[157] = 10'b0101100111;
    16'b0000001110010010: out_v[157] = 10'b1000000110;
    16'b0000001110011000: out_v[157] = 10'b1011100111;
    16'b0000101110010000: out_v[157] = 10'b1101010110;
    16'b0000001000010000: out_v[157] = 10'b1100001011;
    16'b0100001110010000: out_v[157] = 10'b1110100011;
    16'b0000100100011010: out_v[157] = 10'b0000011111;
    16'b0100000110001000: out_v[157] = 10'b1101000110;
    16'b0000001100010010: out_v[157] = 10'b1110110011;
    16'b0000001000010010: out_v[157] = 10'b0111011001;
    16'b0000001010010010: out_v[157] = 10'b1111001010;
    16'b0100101110001000: out_v[157] = 10'b1111010111;
    16'b0100101100001010: out_v[157] = 10'b0110110110;
    16'b0100101010011000: out_v[157] = 10'b1110101010;
    16'b0100100110001000: out_v[157] = 10'b1000101101;
    16'b0000001010000010: out_v[157] = 10'b1010010100;
    16'b0000101010001000: out_v[157] = 10'b0111101010;
    16'b0000001010001000: out_v[157] = 10'b1100001100;
    16'b0100001010011010: out_v[157] = 10'b0101010010;
    16'b0000101010011010: out_v[157] = 10'b1010010011;
    16'b0100001010001000: out_v[157] = 10'b1101010110;
    16'b0000001010011010: out_v[157] = 10'b0100001010;
    16'b0100101010001000: out_v[157] = 10'b1011011010;
    16'b0000001110011010: out_v[157] = 10'b1101101011;
    16'b0100100010001000: out_v[157] = 10'b0001101101;
    16'b0100001000011000: out_v[157] = 10'b1001011101;
    16'b0100001000001000: out_v[157] = 10'b0111011001;
    16'b0000101110011010: out_v[157] = 10'b1010001110;
    16'b0100101000001000: out_v[157] = 10'b0111011010;
    16'b0000101010000000: out_v[157] = 10'b1001110111;
    16'b0000001110001000: out_v[157] = 10'b1011101101;
    16'b0000001010001010: out_v[157] = 10'b0011111101;
    16'b0000101010001010: out_v[157] = 10'b1100001011;
    16'b0000101110001010: out_v[157] = 10'b1000101011;
    16'b0100101010000000: out_v[157] = 10'b0110011111;
    16'b0000101010000010: out_v[157] = 10'b1001001010;
    16'b0100101010001001: out_v[157] = 10'b0100111010;
    16'b0100101010001010: out_v[157] = 10'b0100100010;
    16'b0100101000011000: out_v[157] = 10'b1101000010;
    16'b0000000110001000: out_v[157] = 10'b0010011011;
    16'b0000000000011000: out_v[157] = 10'b0001010011;
    16'b0000000110011010: out_v[157] = 10'b0000010001;
    16'b0000000010001000: out_v[157] = 10'b0011000010;
    16'b0100000100011000: out_v[157] = 10'b1111001010;
    16'b0000100110001000: out_v[157] = 10'b1000111100;
    16'b0000000110010000: out_v[157] = 10'b0011111010;
    16'b0000000110001010: out_v[157] = 10'b1101011000;
    16'b0000000110011000: out_v[157] = 10'b0101011000;
    16'b0000100100001000: out_v[157] = 10'b0011010111;
    16'b0000000000011010: out_v[157] = 10'b0011110111;
    16'b0000000100001000: out_v[157] = 10'b0000011100;
    16'b0000000010011010: out_v[157] = 10'b1101011000;
    16'b0000100100001010: out_v[157] = 10'b0000111011;
    16'b0000000100001010: out_v[157] = 10'b0010011011;
    16'b0000000110010010: out_v[157] = 10'b0011100010;
    16'b0100001110001000: out_v[157] = 10'b0001110010;
    16'b0000000000001010: out_v[157] = 10'b1001111101;
    16'b0000000010011000: out_v[157] = 10'b0001001111;
    16'b0000000100011000: out_v[157] = 10'b0000011101;
    16'b0000000000001000: out_v[157] = 10'b0001110010;
    16'b0000000000010010: out_v[157] = 10'b1000010111;
    16'b0100000110011000: out_v[157] = 10'b1111100001;
    16'b0100000110001010: out_v[157] = 10'b1000011101;
    16'b0000000100010010: out_v[157] = 10'b0111011111;
    16'b0000000110000000: out_v[157] = 10'b0000110111;
    16'b0000100110001010: out_v[157] = 10'b0110010001;
    16'b0100000010011000: out_v[157] = 10'b1001100010;
    16'b0100000000010010: out_v[157] = 10'b1001101101;
    16'b0100000110010000: out_v[157] = 10'b0110001101;
    16'b0100001000010010: out_v[157] = 10'b0001111100;
    16'b0000101000001000: out_v[157] = 10'b1010100000;
    16'b0100000100010010: out_v[157] = 10'b1100101100;
    16'b0100000010010010: out_v[157] = 10'b0110000101;
    16'b0100000110010010: out_v[157] = 10'b1001101100;
    16'b0100001100010010: out_v[157] = 10'b0000110011;
    16'b0100001000001010: out_v[157] = 10'b1101010010;
    16'b0000001000001000: out_v[157] = 10'b0000100110;
    16'b0100001100000010: out_v[157] = 10'b1101101110;
    16'b0100101000001010: out_v[157] = 10'b1001110010;
    16'b0100000100000010: out_v[157] = 10'b1101101000;
    16'b0000101000001010: out_v[157] = 10'b1100100010;
    16'b0100000000011000: out_v[157] = 10'b0111110110;
    16'b0000001000001010: out_v[157] = 10'b1001001110;
    16'b0100000010011010: out_v[157] = 10'b0000000110;
    16'b0100000000000010: out_v[157] = 10'b1101100001;
    16'b0000100110011000: out_v[157] = 10'b1011001010;
    16'b0000100100011000: out_v[157] = 10'b1011101110;
    16'b0000100000011000: out_v[157] = 10'b0101010000;
    16'b0000100010010000: out_v[157] = 10'b1111100010;
    16'b0000100000010000: out_v[157] = 10'b1011001010;
    16'b0000100100010000: out_v[157] = 10'b1101100011;
    16'b0000100110010000: out_v[157] = 10'b0001000010;
    16'b0000000100010000: out_v[157] = 10'b0011101001;
    16'b0100001100010000: out_v[157] = 10'b0001010101;
    16'b0100000010001000: out_v[157] = 10'b1001000111;
    16'b0100001010000010: out_v[157] = 10'b1011111000;
    16'b0100100010011000: out_v[157] = 10'b0110011000;
    16'b0100000000001000: out_v[157] = 10'b1110101011;
    16'b0100000100001000: out_v[157] = 10'b1011001110;
    16'b0100001110010010: out_v[157] = 10'b1100010111;
    16'b0100001110001010: out_v[157] = 10'b1101000011;
    16'b0000001110000010: out_v[157] = 10'b0111010000;
    16'b0100001010001010: out_v[157] = 10'b0100110101;
    16'b0100001110000000: out_v[157] = 10'b0100111100;
    16'b0100001110000010: out_v[157] = 10'b0111010110;
    16'b0000001110001010: out_v[157] = 10'b1010001101;
    16'b0100000110000000: out_v[157] = 10'b1100001100;
    default: out_v[157] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000001010100000: out_v[158] = 10'b1001001000;
    16'b0000001100101000: out_v[158] = 10'b1001000011;
    16'b0000001110001000: out_v[158] = 10'b1100111111;
    16'b0000001110111000: out_v[158] = 10'b1011001011;
    16'b0000000010001000: out_v[158] = 10'b0111110110;
    16'b0000001000000000: out_v[158] = 10'b1010101101;
    16'b0000001111001000: out_v[158] = 10'b0010001011;
    16'b0000001100001000: out_v[158] = 10'b1011011100;
    16'b0000001000111000: out_v[158] = 10'b1101110100;
    16'b0000001000100000: out_v[158] = 10'b1000011111;
    16'b0000001100111000: out_v[158] = 10'b0011110000;
    16'b0000001000101000: out_v[158] = 10'b0010111001;
    16'b0000001100110000: out_v[158] = 10'b1101011010;
    16'b0000001110101000: out_v[158] = 10'b0010101111;
    16'b0000001010101000: out_v[158] = 10'b0000110011;
    16'b0000001010001000: out_v[158] = 10'b1010100000;
    16'b0000001000001000: out_v[158] = 10'b1101011111;
    16'b0000001110100000: out_v[158] = 10'b1111000111;
    16'b0000000110101000: out_v[158] = 10'b0010101110;
    16'b0000001111101000: out_v[158] = 10'b1001110000;
    16'b0000001100100000: out_v[158] = 10'b1100110111;
    16'b0000001100000000: out_v[158] = 10'b0000011011;
    16'b0000001010111000: out_v[158] = 10'b0000100101;
    16'b0000000110011000: out_v[158] = 10'b0000001011;
    16'b0000000110001000: out_v[158] = 10'b1100010001;
    16'b0000000100001000: out_v[158] = 10'b1001010111;
    16'b0000001111100000: out_v[158] = 10'b1100010101;
    16'b0000001000110000: out_v[158] = 10'b0001000011;
    16'b0010000000000000: out_v[158] = 10'b0111111011;
    16'b0010001000100000: out_v[158] = 10'b1111001010;
    16'b0010001000000000: out_v[158] = 10'b1100011010;
    16'b0010000000010000: out_v[158] = 10'b1110101101;
    16'b0010001000010000: out_v[158] = 10'b1011101010;
    16'b0010000010000000: out_v[158] = 10'b0001010111;
    16'b0010001010100000: out_v[158] = 10'b0100001101;
    16'b0010001000110000: out_v[158] = 10'b1011010110;
    16'b0000000000000000: out_v[158] = 10'b0001111110;
    16'b0010000100000000: out_v[158] = 10'b0011010110;
    16'b0010000100110000: out_v[158] = 10'b1011101011;
    16'b0010001100110000: out_v[158] = 10'b1001000111;
    16'b0010001010000000: out_v[158] = 10'b0110100100;
    16'b0010000100010000: out_v[158] = 10'b1110101001;
    16'b0000000000010000: out_v[158] = 10'b1110010110;
    16'b0010001100100000: out_v[158] = 10'b0100011110;
    16'b0010000110010000: out_v[158] = 10'b0011001111;
    16'b0010001110101000: out_v[158] = 10'b0110000110;
    16'b0010001010110000: out_v[158] = 10'b0110000110;
    16'b0010000100011000: out_v[158] = 10'b1100101100;
    16'b0010001100101000: out_v[158] = 10'b1100111110;
    16'b0010101110100000: out_v[158] = 10'b1010111100;
    16'b0010001110110000: out_v[158] = 10'b0111011110;
    16'b0010001100000000: out_v[158] = 10'b1111011010;
    16'b0010001100111000: out_v[158] = 10'b1011110011;
    16'b0010001110100000: out_v[158] = 10'b1000000100;
    16'b0010000000100000: out_v[158] = 10'b0111001000;
    16'b0010000000110000: out_v[158] = 10'b1100100101;
    16'b0000000100010000: out_v[158] = 10'b1010011100;
    16'b0010000010010000: out_v[158] = 10'b1111011000;
    16'b0010000010110000: out_v[158] = 10'b0001001010;
    16'b0010101010100000: out_v[158] = 10'b1111110111;
    16'b0010001110111000: out_v[158] = 10'b0001011011;
    16'b0010001000101000: out_v[158] = 10'b0000111111;
    16'b0010001110000000: out_v[158] = 10'b0101110111;
    16'b0000000000110000: out_v[158] = 10'b1001111000;
    16'b0000000000001000: out_v[158] = 10'b1101001011;
    16'b0010001010101000: out_v[158] = 10'b1100101001;
    16'b0000000010100000: out_v[158] = 10'b1111000011;
    16'b0000001010000000: out_v[158] = 10'b0011100001;
    16'b0000000000100000: out_v[158] = 10'b1001011010;
    16'b0000001010110000: out_v[158] = 10'b1001010111;
    16'b0000000000011000: out_v[158] = 10'b0010110100;
    16'b0010000010001000: out_v[158] = 10'b0000010010;
    16'b0000000010000000: out_v[158] = 10'b0000110010;
    16'b0010000000001000: out_v[158] = 10'b1101110100;
    16'b0010000110001000: out_v[158] = 10'b0001111000;
    16'b0010000100001000: out_v[158] = 10'b1101011010;
    16'b0010001010001000: out_v[158] = 10'b1110000101;
    16'b0010000110000000: out_v[158] = 10'b0100010110;
    16'b0010001000001000: out_v[158] = 10'b0001110000;
    16'b0000000100000000: out_v[158] = 10'b0101100011;
    16'b0000001110000000: out_v[158] = 10'b0010111110;
    16'b0000000010010000: out_v[158] = 10'b1101100111;
    16'b0000000010011000: out_v[158] = 10'b0011101010;
    16'b0000000010110000: out_v[158] = 10'b1100110111;
    16'b0010001000111000: out_v[158] = 10'b1111100001;
    16'b0000001000010000: out_v[158] = 10'b0100100100;
    16'b0010000011001000: out_v[158] = 10'b0001111001;
    16'b0010001010111000: out_v[158] = 10'b1011011000;
    16'b0010000010011000: out_v[158] = 10'b1001001111;
    16'b0010001100001000: out_v[158] = 10'b1101001110;
    16'b0000000010000001: out_v[158] = 10'b0101011000;
    16'b0000001010000001: out_v[158] = 10'b0111010111;
    16'b0000000000000001: out_v[158] = 10'b0010111111;
    16'b0000000000001101: out_v[158] = 10'b0011000110;
    16'b0000000000000101: out_v[158] = 10'b0001110111;
    16'b0000001010001001: out_v[158] = 10'b1001101001;
    16'b0000000000001001: out_v[158] = 10'b1011011001;
    16'b0000000010001001: out_v[158] = 10'b0100011000;
    16'b0010000010100000: out_v[158] = 10'b1100000111;
    default: out_v[158] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001000100100000: out_v[159] = 10'b1001100111;
    16'b0001000000100000: out_v[159] = 10'b0001010011;
    16'b0001000100110010: out_v[159] = 10'b0011011000;
    16'b1000000100100010: out_v[159] = 10'b1100011111;
    16'b0001000000100010: out_v[159] = 10'b1001000001;
    16'b0000000000100000: out_v[159] = 10'b1000111011;
    16'b0001010000100010: out_v[159] = 10'b0000000111;
    16'b0000000000000010: out_v[159] = 10'b0110100111;
    16'b0000000000100010: out_v[159] = 10'b0101110111;
    16'b0001000100100010: out_v[159] = 10'b1001010011;
    16'b1000000000000000: out_v[159] = 10'b0010010111;
    16'b0001000000110010: out_v[159] = 10'b0101011100;
    16'b0001010000110000: out_v[159] = 10'b0111000011;
    16'b1000000000100000: out_v[159] = 10'b1000110011;
    16'b0000000100100010: out_v[159] = 10'b1100100011;
    16'b0000000000110000: out_v[159] = 10'b1000101000;
    16'b1001000000100000: out_v[159] = 10'b1001010101;
    16'b0001010100100010: out_v[159] = 10'b0011010011;
    16'b0001000000110000: out_v[159] = 10'b0011101101;
    16'b0000000000000000: out_v[159] = 10'b0110010010;
    16'b1001000000110000: out_v[159] = 10'b0111011000;
    16'b1000000000100010: out_v[159] = 10'b1011010111;
    16'b0000000000000011: out_v[159] = 10'b0011110111;
    16'b1000000000000010: out_v[159] = 10'b1101010010;
    16'b0101001100100010: out_v[159] = 10'b1110001011;
    16'b0001000000000000: out_v[159] = 10'b1111001010;
    16'b1001000000100010: out_v[159] = 10'b1111010111;
    16'b0000000100000010: out_v[159] = 10'b0010011001;
    16'b0000000100110010: out_v[159] = 10'b1010001001;
    16'b0000000000110010: out_v[159] = 10'b0101101001;
    16'b0001010000100000: out_v[159] = 10'b0100010100;
    16'b1001000100100010: out_v[159] = 10'b1000110111;
    16'b0001010000110010: out_v[159] = 10'b1001010111;
    16'b1001010000110000: out_v[159] = 10'b0011001011;
    16'b0000010000010000: out_v[159] = 10'b0111100001;
    16'b0000000000010000: out_v[159] = 10'b1000001100;
    16'b1000010000110000: out_v[159] = 10'b0110010111;
    16'b0000010000110000: out_v[159] = 10'b1101010011;
    16'b0000000100010000: out_v[159] = 10'b1000010011;
    16'b0000010100010000: out_v[159] = 10'b0101000111;
    16'b1000010000010000: out_v[159] = 10'b1001010101;
    16'b0001010000110001: out_v[159] = 10'b0110110010;
    16'b0000010100110000: out_v[159] = 10'b1011010111;
    16'b0001010100110000: out_v[159] = 10'b0110100101;
    16'b0001010100100000: out_v[159] = 10'b0011010010;
    16'b1001010000100000: out_v[159] = 10'b1111000110;
    16'b0101011000110000: out_v[159] = 10'b1010001010;
    16'b0000010100100000: out_v[159] = 10'b1010110100;
    16'b0000000100000000: out_v[159] = 10'b0111000101;
    16'b1001010000100001: out_v[159] = 10'b1000110100;
    16'b0000010000100000: out_v[159] = 10'b0100110101;
    16'b0000010000100010: out_v[159] = 10'b1000101111;
    16'b1001010100100000: out_v[159] = 10'b1001010100;
    16'b0000010000000000: out_v[159] = 10'b1101001001;
    16'b0101011100110000: out_v[159] = 10'b1001110110;
    16'b0101011000100000: out_v[159] = 10'b0011011010;
    16'b0100011000100000: out_v[159] = 10'b1111011000;
    16'b0101011000110010: out_v[159] = 10'b0111111010;
    16'b1001010100110000: out_v[159] = 10'b1001000111;
    16'b0000010100000000: out_v[159] = 10'b1101101111;
    16'b1000010100100000: out_v[159] = 10'b1010101100;
    16'b0000000100100000: out_v[159] = 10'b1001111110;
    16'b0101011000100010: out_v[159] = 10'b1001111001;
    16'b0001010000010010: out_v[159] = 10'b0110110111;
    16'b0001010000000000: out_v[159] = 10'b1000111000;
    16'b0001010000000010: out_v[159] = 10'b0111001011;
    16'b1000010000100000: out_v[159] = 10'b1110100010;
    16'b0001010100000000: out_v[159] = 10'b0000101000;
    16'b1001010100100001: out_v[159] = 10'b0111110011;
    16'b1001010000100010: out_v[159] = 10'b1101000001;
    16'b0001010000100001: out_v[159] = 10'b1010000110;
    16'b0000000100010001: out_v[159] = 10'b1000100001;
    16'b0000000100110000: out_v[159] = 10'b1001001011;
    16'b0000000000010001: out_v[159] = 10'b0001001101;
    16'b0001000100110000: out_v[159] = 10'b0100101010;
    16'b0000000100010010: out_v[159] = 10'b0000111100;
    16'b1000000000010001: out_v[159] = 10'b1101001100;
    16'b1000000000110000: out_v[159] = 10'b0010100000;
    16'b1000000000110001: out_v[159] = 10'b1111010100;
    16'b0000000000110001: out_v[159] = 10'b1001011110;
    16'b0000000100010011: out_v[159] = 10'b0101001111;
    16'b0000000000010010: out_v[159] = 10'b1110011110;
    16'b1000000000010000: out_v[159] = 10'b1100100100;
    16'b0001010100000010: out_v[159] = 10'b0100110010;
    16'b1000010000000000: out_v[159] = 10'b1001011111;
    16'b0000010000010010: out_v[159] = 10'b1000010100;
    16'b0000010000000010: out_v[159] = 10'b0111100011;
    16'b1001010000000000: out_v[159] = 10'b1010110110;
    16'b0001010000010000: out_v[159] = 10'b1000111000;
    16'b1001010100000000: out_v[159] = 10'b0010110010;
    16'b1001000100110000: out_v[159] = 10'b1110110001;
    16'b0000000000000001: out_v[159] = 10'b1011110000;
    16'b1000000100110000: out_v[159] = 10'b0010010111;
    16'b1000000100110010: out_v[159] = 10'b1010111110;
    16'b1001010100100010: out_v[159] = 10'b0111010011;
    16'b0001010100110010: out_v[159] = 10'b0111010000;
    16'b0001000000000010: out_v[159] = 10'b0101100000;
    16'b1001010000010000: out_v[159] = 10'b0100001010;
    16'b1001010000110010: out_v[159] = 10'b0101101101;
    16'b0001010100010000: out_v[159] = 10'b0001101101;
    16'b0000010000100001: out_v[159] = 10'b1011100001;
    16'b0001010000010001: out_v[159] = 10'b1101011010;
    16'b0001000100010000: out_v[159] = 10'b1110000110;
    16'b0001000000010000: out_v[159] = 10'b0110101110;
    default: out_v[159] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001000100000011: out_v[160] = 10'b1001100111;
    16'b0001000001100001: out_v[160] = 10'b1110011101;
    16'b0001000100001011: out_v[160] = 10'b1011011001;
    16'b0001000010000001: out_v[160] = 10'b1101010000;
    16'b0000101000000010: out_v[160] = 10'b1011010111;
    16'b0000101001101010: out_v[160] = 10'b0011101000;
    16'b0001000110001011: out_v[160] = 10'b1011001011;
    16'b0001000000100001: out_v[160] = 10'b0101011001;
    16'b0001001001100001: out_v[160] = 10'b1110100011;
    16'b0001100001100011: out_v[160] = 10'b0111010111;
    16'b0000000001100011: out_v[160] = 10'b0010110110;
    16'b0001000000000010: out_v[160] = 10'b1010000101;
    16'b0001100000000010: out_v[160] = 10'b1001011000;
    16'b0001000000001011: out_v[160] = 10'b0001100001;
    16'b0001000000100011: out_v[160] = 10'b1101010011;
    16'b0001000000000011: out_v[160] = 10'b1011101011;
    16'b0001000000101011: out_v[160] = 10'b1110111011;
    16'b0000101001100010: out_v[160] = 10'b0111011011;
    16'b0001101001100010: out_v[160] = 10'b1000111111;
    16'b0001101001101010: out_v[160] = 10'b1101110011;
    16'b0001000000001001: out_v[160] = 10'b1110100001;
    16'b0000000001100001: out_v[160] = 10'b0010011111;
    16'b0001101001100011: out_v[160] = 10'b1110011011;
    16'b0001100000001010: out_v[160] = 10'b0111111111;
    16'b0000000000001011: out_v[160] = 10'b0010100011;
    16'b0000100000001000: out_v[160] = 10'b1111111101;
    16'b0001000000000001: out_v[160] = 10'b1001011001;
    16'b0000100001100010: out_v[160] = 10'b1111001110;
    16'b0000100000000010: out_v[160] = 10'b0010111000;
    16'b0000101001100011: out_v[160] = 10'b0110000111;
    16'b0001000000001010: out_v[160] = 10'b0111110010;
    16'b0001000001101011: out_v[160] = 10'b1001101011;
    16'b0001000000001000: out_v[160] = 10'b0011011000;
    16'b0000100001100011: out_v[160] = 10'b1000011110;
    16'b0001000001100011: out_v[160] = 10'b1011011011;
    16'b0001000010001011: out_v[160] = 10'b0011000001;
    16'b0000101000001010: out_v[160] = 10'b1101010011;
    16'b0000100001101010: out_v[160] = 10'b1111001110;
    16'b0001000110000011: out_v[160] = 10'b0010111101;
    16'b0000101001000010: out_v[160] = 10'b1111111110;
    16'b0000000000001010: out_v[160] = 10'b1000011010;
    16'b0000101001100000: out_v[160] = 10'b1001011111;
    16'b0000100000001010: out_v[160] = 10'b1011011010;
    16'b0001101001101011: out_v[160] = 10'b1111101111;
    16'b0000000110000000: out_v[160] = 10'b1001010011;
    16'b0000000000000000: out_v[160] = 10'b1100100111;
    16'b0000000000000010: out_v[160] = 10'b0001111001;
    16'b0000000000001000: out_v[160] = 10'b0100001011;
    16'b0000000100000000: out_v[160] = 10'b0010001011;
    16'b0100000000000010: out_v[160] = 10'b0111110101;
    16'b0000000000000001: out_v[160] = 10'b1011001110;
    16'b0000000100000001: out_v[160] = 10'b1111001100;
    16'b0000000100001010: out_v[160] = 10'b1110010001;
    16'b0000000100001000: out_v[160] = 10'b1100111101;
    16'b0000000110100000: out_v[160] = 10'b1110011111;
    16'b0000000010001000: out_v[160] = 10'b0000011010;
    16'b0000000110001000: out_v[160] = 10'b1100010110;
    16'b0000000110000001: out_v[160] = 10'b1001101011;
    16'b0000000010000000: out_v[160] = 10'b1110000010;
    16'b0000000000000011: out_v[160] = 10'b0110101011;
    16'b0100000110000010: out_v[160] = 10'b1011111111;
    16'b0100000110001010: out_v[160] = 10'b1101110001;
    16'b0101000010001001: out_v[160] = 10'b1110100101;
    16'b0100000110001000: out_v[160] = 10'b1010101100;
    16'b0100000100001000: out_v[160] = 10'b1100110101;
    16'b0101000110001000: out_v[160] = 10'b1111010111;
    16'b0000000010000010: out_v[160] = 10'b1000011101;
    16'b0001000110000000: out_v[160] = 10'b1101000101;
    16'b0100000110000000: out_v[160] = 10'b1000110111;
    16'b0000000110001010: out_v[160] = 10'b0010111101;
    16'b0000000110100010: out_v[160] = 10'b1011010100;
    16'b0100000010001000: out_v[160] = 10'b1110010101;
    16'b0101000100001000: out_v[160] = 10'b0100000100;
    16'b0001000110000010: out_v[160] = 10'b0010100111;
    16'b0101000110001010: out_v[160] = 10'b1111011010;
    16'b0001000110001000: out_v[160] = 10'b0001001100;
    16'b0001000100001010: out_v[160] = 10'b1001111110;
    16'b0000000100000010: out_v[160] = 10'b0111110100;
    16'b0101000010001000: out_v[160] = 10'b1111100111;
    16'b0000000100001011: out_v[160] = 10'b1011010010;
    16'b0001000110001010: out_v[160] = 10'b1100010010;
    16'b0001000100000010: out_v[160] = 10'b0010100100;
    16'b0000000110000010: out_v[160] = 10'b1001000110;
    16'b0000000100000011: out_v[160] = 10'b1110011000;
    16'b0100000100001001: out_v[160] = 10'b0100100110;
    16'b0000000010001010: out_v[160] = 10'b0001111110;
    16'b0000000110001011: out_v[160] = 10'b0011010011;
    16'b0000100110000010: out_v[160] = 10'b1001001110;
    16'b0101000000001000: out_v[160] = 10'b1010100110;
    16'b0100000010001001: out_v[160] = 10'b0011011111;
    16'b0001000010000011: out_v[160] = 10'b0010011110;
    16'b0000000000000111: out_v[160] = 10'b1011101000;
    16'b0001000010110011: out_v[160] = 10'b1100100011;
    16'b0000000110000011: out_v[160] = 10'b1001011011;
    16'b0001000000000111: out_v[160] = 10'b0010011011;
    16'b0001000010000111: out_v[160] = 10'b1000011110;
    16'b0000000010001011: out_v[160] = 10'b1101110100;
    16'b0001000010001001: out_v[160] = 10'b0100101001;
    16'b0101000010001011: out_v[160] = 10'b1110111001;
    16'b0001000010100011: out_v[160] = 10'b0011110110;
    16'b0001000010000010: out_v[160] = 10'b0011110001;
    16'b0000000010000011: out_v[160] = 10'b0010101100;
    16'b0001000010000000: out_v[160] = 10'b0100111001;
    16'b0100000000001001: out_v[160] = 10'b1010001111;
    16'b0001000010001000: out_v[160] = 10'b1001001100;
    16'b0101000010000011: out_v[160] = 10'b0010011001;
    16'b0101000010000001: out_v[160] = 10'b0101100111;
    16'b0101000000001001: out_v[160] = 10'b1110011110;
    16'b0000000000001001: out_v[160] = 10'b1100011100;
    16'b0001000010001010: out_v[160] = 10'b1001110001;
    16'b0000000010001001: out_v[160] = 10'b0100101010;
    16'b0001000010010011: out_v[160] = 10'b0111111010;
    16'b0000000010000001: out_v[160] = 10'b0010111101;
    16'b0001100010000011: out_v[160] = 10'b1001001101;
    16'b0001100110000101: out_v[160] = 10'b1100010101;
    16'b0001000110000001: out_v[160] = 10'b0101000010;
    16'b0001000100000001: out_v[160] = 10'b0010111110;
    16'b0000000010100001: out_v[160] = 10'b1111000011;
    16'b0001100010000100: out_v[160] = 10'b1000011010;
    16'b0000100010000101: out_v[160] = 10'b1101010011;
    16'b0001101110000000: out_v[160] = 10'b0000110001;
    16'b0001100010000101: out_v[160] = 10'b0011011011;
    16'b0001000110100011: out_v[160] = 10'b0100100011;
    16'b0001100110000001: out_v[160] = 10'b0111100111;
    16'b0001100110100000: out_v[160] = 10'b0110110011;
    16'b0001100010000001: out_v[160] = 10'b0010110111;
    16'b0001101010100001: out_v[160] = 10'b1001011111;
    16'b0000100110000100: out_v[160] = 10'b1101101110;
    16'b0001100110000000: out_v[160] = 10'b0100100111;
    16'b0001100010000000: out_v[160] = 10'b1101110011;
    16'b0001000010100001: out_v[160] = 10'b0100110110;
    16'b0001100110000100: out_v[160] = 10'b0111101111;
    16'b0001000110000101: out_v[160] = 10'b0100110010;
    16'b0000100010000001: out_v[160] = 10'b0010011001;
    16'b0001000110100001: out_v[160] = 10'b1001100111;
    16'b0001101110000100: out_v[160] = 10'b1010111111;
    16'b0000000110100001: out_v[160] = 10'b0100010010;
    16'b0000100110000000: out_v[160] = 10'b0001001110;
    16'b0000000010000101: out_v[160] = 10'b0101010111;
    16'b0001101010000001: out_v[160] = 10'b0110001011;
    16'b0001101010000101: out_v[160] = 10'b1000111101;
    16'b0001101010000000: out_v[160] = 10'b1001100001;
    16'b0001101110100000: out_v[160] = 10'b0110111111;
    16'b0000000001000001: out_v[160] = 10'b0010110010;
    16'b0000000000100001: out_v[160] = 10'b0100100100;
    16'b0000000000100011: out_v[160] = 10'b1101010110;
    16'b0000000101100001: out_v[160] = 10'b1011101000;
    16'b0001100010100011: out_v[160] = 10'b0101101110;
    16'b0000000100100001: out_v[160] = 10'b1001101000;
    16'b0000000000100000: out_v[160] = 10'b0111100001;
    16'b0000000100100011: out_v[160] = 10'b1100101110;
    16'b0001100010000111: out_v[160] = 10'b1100100111;
    16'b0000100000100001: out_v[160] = 10'b0000100010;
    16'b0000100000100011: out_v[160] = 10'b1010010101;
    16'b0000000010100011: out_v[160] = 10'b0010101011;
    16'b0000100000000011: out_v[160] = 10'b1000111001;
    16'b0001100010001011: out_v[160] = 10'b0100110001;
    16'b0101000110001011: out_v[160] = 10'b1001010101;
    16'b0000000100001001: out_v[160] = 10'b0110011101;
    16'b0101000110000011: out_v[160] = 10'b1011110011;
    16'b0001000100001001: out_v[160] = 10'b1110110101;
    16'b0101000110000001: out_v[160] = 10'b1111010011;
    16'b0101100110001000: out_v[160] = 10'b0011010110;
    16'b0001000110001001: out_v[160] = 10'b0100110011;
    16'b0000000110001001: out_v[160] = 10'b1011110011;
    16'b0101000110000000: out_v[160] = 10'b1110101110;
    16'b0100100110000000: out_v[160] = 10'b1110111110;
    16'b0101100110000000: out_v[160] = 10'b0010101010;
    16'b0001100011100000: out_v[160] = 10'b1011101001;
    16'b0001100000000000: out_v[160] = 10'b0101010110;
    16'b0000100010000000: out_v[160] = 10'b0110100100;
    16'b0001000010000100: out_v[160] = 10'b0111110011;
    16'b0001100010000010: out_v[160] = 10'b0010110111;
    16'b0000100010000010: out_v[160] = 10'b1001100100;
    16'b0001100000000100: out_v[160] = 10'b0111001111;
    16'b0001100010000110: out_v[160] = 10'b0010001011;
    16'b0000100010100000: out_v[160] = 10'b0011110011;
    16'b0000000010100000: out_v[160] = 10'b1111000011;
    16'b0000100010000100: out_v[160] = 10'b0010111101;
    16'b0001000010100010: out_v[160] = 10'b0011011011;
    16'b0000000010100010: out_v[160] = 10'b1000011101;
    16'b0001000000000000: out_v[160] = 10'b1100110110;
    16'b0001100010100010: out_v[160] = 10'b0001111011;
    16'b0001100010100000: out_v[160] = 10'b0111100111;
    16'b0001000111100011: out_v[160] = 10'b0100011100;
    16'b0000000111100011: out_v[160] = 10'b0001101110;
    16'b0000000110100011: out_v[160] = 10'b0000010011;
    16'b0000100110100011: out_v[160] = 10'b0111110010;
    16'b0000000111100010: out_v[160] = 10'b0101110011;
    16'b0000000111000011: out_v[160] = 10'b0111010011;
    16'b0000000111100001: out_v[160] = 10'b1101100000;
    16'b0000100010000111: out_v[160] = 10'b1101101001;
    16'b0000100110000011: out_v[160] = 10'b0110100010;
    16'b0000000110000111: out_v[160] = 10'b1000001101;
    16'b0000100111100011: out_v[160] = 10'b0110010111;
    16'b0001100110000111: out_v[160] = 10'b1010000011;
    16'b0000000110101011: out_v[160] = 10'b1100110111;
    16'b0001100110000011: out_v[160] = 10'b0011101010;
    16'b0000100110000111: out_v[160] = 10'b1111110010;
    16'b0000000110000110: out_v[160] = 10'b1011101011;
    16'b0001101110000010: out_v[160] = 10'b0100110010;
    16'b0001101110000110: out_v[160] = 10'b1101110000;
    16'b0001100110000110: out_v[160] = 10'b1001000101;
    16'b0000100010000011: out_v[160] = 10'b1101000111;
    16'b0000000010000111: out_v[160] = 10'b0111000100;
    16'b0000100110000110: out_v[160] = 10'b0000100111;
    16'b0000100010000110: out_v[160] = 10'b1011101100;
    16'b0001100110000010: out_v[160] = 10'b1001000111;
    16'b0000000010000110: out_v[160] = 10'b0000000101;
    16'b0001000110000110: out_v[160] = 10'b0111111010;
    default: out_v[160] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010000000000000: out_v[161] = 10'b0111011101;
    16'b0110010000000100: out_v[161] = 10'b1001101111;
    16'b0100010000000000: out_v[161] = 10'b0110110101;
    16'b0010010000000000: out_v[161] = 10'b1001110010;
    16'b0010010000000001: out_v[161] = 10'b1000101010;
    16'b0110010000000001: out_v[161] = 10'b0001000011;
    16'b0110010000000000: out_v[161] = 10'b0101000010;
    16'b0000010000000000: out_v[161] = 10'b1110111101;
    16'b0100010000000100: out_v[161] = 10'b1101000011;
    16'b0010010000000100: out_v[161] = 10'b0110000111;
    16'b0100010000000001: out_v[161] = 10'b0010010110;
    16'b0000010000000100: out_v[161] = 10'b0101111001;
    16'b0110010000100000: out_v[161] = 10'b1011011111;
    16'b0010000000000001: out_v[161] = 10'b0011011100;
    16'b0100000000000000: out_v[161] = 10'b0000111101;
    16'b0100110000000000: out_v[161] = 10'b0111011101;
    16'b0110110000000000: out_v[161] = 10'b1010010011;
    16'b0000010000000001: out_v[161] = 10'b0101000110;
    16'b0010000000000100: out_v[161] = 10'b0111000101;
    16'b0000000000000000: out_v[161] = 10'b1000111000;
    16'b0110110000100000: out_v[161] = 10'b0010010001;
    16'b0010110000000000: out_v[161] = 10'b0011110100;
    16'b0000000000000101: out_v[161] = 10'b1011110011;
    16'b0000000000000001: out_v[161] = 10'b0111010111;
    16'b0010000000000101: out_v[161] = 10'b1001101110;
    16'b0000000000000100: out_v[161] = 10'b0001101100;
    16'b0010100000000000: out_v[161] = 10'b0110110100;
    16'b0000100000000001: out_v[161] = 10'b1101010110;
    16'b0010110000001001: out_v[161] = 10'b0101000011;
    16'b0000000000100001: out_v[161] = 10'b1110000111;
    16'b0010110000100001: out_v[161] = 10'b1011011111;
    16'b0010000000100001: out_v[161] = 10'b0000111110;
    16'b0010110000000001: out_v[161] = 10'b1010001000;
    16'b0000110000000001: out_v[161] = 10'b0111010111;
    16'b0010100000000001: out_v[161] = 10'b0011000100;
    16'b0010010000001001: out_v[161] = 10'b1010111111;
    16'b0000100000100001: out_v[161] = 10'b0100000101;
    16'b0000100000000000: out_v[161] = 10'b1010111010;
    16'b0000110000000000: out_v[161] = 10'b1111101100;
    16'b0010100000100001: out_v[161] = 10'b0000110111;
    16'b0000000000100100: out_v[161] = 10'b0000011111;
    16'b0000000000100000: out_v[161] = 10'b1010000010;
    16'b0000100000100000: out_v[161] = 10'b1011110000;
    16'b0010000000100000: out_v[161] = 10'b1010011011;
    16'b0000010000000101: out_v[161] = 10'b0111010010;
    16'b0100000000000001: out_v[161] = 10'b0110011010;
    16'b0110000000000001: out_v[161] = 10'b0011100100;
    16'b0111010000000001: out_v[161] = 10'b0110101111;
    16'b0000000000100101: out_v[161] = 10'b0110110011;
    16'b0000000010100000: out_v[161] = 10'b1110010111;
    16'b0000000010000000: out_v[161] = 10'b1001001010;
    16'b0010010000000101: out_v[161] = 10'b1100110000;
    16'b0110000000000000: out_v[161] = 10'b0101001010;
    16'b0010100000100000: out_v[161] = 10'b1100010011;
    default: out_v[161] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010000000000010: out_v[162] = 10'b1001010110;
    16'b0011100100000010: out_v[162] = 10'b1011001011;
    16'b0010000000000001: out_v[162] = 10'b0110101011;
    16'b0010000000000011: out_v[162] = 10'b1011100111;
    16'b0000000000000000: out_v[162] = 10'b0010100111;
    16'b0001000000000010: out_v[162] = 10'b1010011011;
    16'b0001000000000000: out_v[162] = 10'b1010100001;
    16'b0011000000000000: out_v[162] = 10'b1100100011;
    16'b0011000000000001: out_v[162] = 10'b0011010001;
    16'b0011000000000010: out_v[162] = 10'b0100100111;
    16'b0010000001000010: out_v[162] = 10'b0101111101;
    16'b0011000100000000: out_v[162] = 10'b1011011110;
    16'b0010000100000010: out_v[162] = 10'b1001010111;
    16'b0010000000000000: out_v[162] = 10'b0111001101;
    16'b0000000000000010: out_v[162] = 10'b0110010101;
    16'b0010100100000010: out_v[162] = 10'b0000101111;
    16'b0010000100000011: out_v[162] = 10'b0101100101;
    16'b0000000000000001: out_v[162] = 10'b0001101000;
    16'b0010000100000000: out_v[162] = 10'b0111000100;
    16'b0011000000000011: out_v[162] = 10'b0000111101;
    16'b0001000000000001: out_v[162] = 10'b1100010011;
    16'b0011000100000001: out_v[162] = 10'b1001101111;
    16'b0000000000000011: out_v[162] = 10'b1011011111;
    16'b0011100100000000: out_v[162] = 10'b0001110011;
    16'b0010000100000001: out_v[162] = 10'b0001110110;
    16'b0011000100000010: out_v[162] = 10'b0011011100;
    16'b0011000001000010: out_v[162] = 10'b1111100101;
    16'b0000000001000000: out_v[162] = 10'b1000011100;
    16'b0000000101000000: out_v[162] = 10'b1010111000;
    16'b0000100000000000: out_v[162] = 10'b0001110111;
    16'b0010000101000000: out_v[162] = 10'b1100000110;
    16'b0010000001000000: out_v[162] = 10'b1100000110;
    16'b0000100101000000: out_v[162] = 10'b0111100100;
    16'b0000100001000000: out_v[162] = 10'b0010100110;
    16'b0000000100000000: out_v[162] = 10'b1001100010;
    16'b0000000001010001: out_v[162] = 10'b1001000111;
    16'b0010000001010000: out_v[162] = 10'b1001001111;
    16'b0000000001000001: out_v[162] = 10'b1110011100;
    16'b0010000001010001: out_v[162] = 10'b0111001000;
    16'b0010000001000001: out_v[162] = 10'b0111010111;
    16'b0000000001000010: out_v[162] = 10'b0101111000;
    16'b0000000001010011: out_v[162] = 10'b1111110100;
    16'b0010000001000011: out_v[162] = 10'b0100111000;
    16'b0010000000010010: out_v[162] = 10'b1010101110;
    16'b0010000001010011: out_v[162] = 10'b1101110010;
    16'b0000000001000011: out_v[162] = 10'b0010100100;
    16'b0010000001110000: out_v[162] = 10'b0001110110;
    16'b0010001001000001: out_v[162] = 10'b1110010101;
    16'b0010000000010011: out_v[162] = 10'b1001100101;
    16'b0010000101000001: out_v[162] = 10'b0001111100;
    16'b0010000101000011: out_v[162] = 10'b0101011000;
    16'b0010000001010010: out_v[162] = 10'b1111001101;
    16'b0000000101010001: out_v[162] = 10'b0001111100;
    16'b0010000101010011: out_v[162] = 10'b1100101110;
    16'b0010100101000011: out_v[162] = 10'b1111011111;
    16'b0000000101000011: out_v[162] = 10'b0011100000;
    16'b0000000101010011: out_v[162] = 10'b1111010010;
    16'b0000000101000001: out_v[162] = 10'b0110101011;
    16'b0000100101000011: out_v[162] = 10'b1100111000;
    16'b0000100101000001: out_v[162] = 10'b0100010110;
    16'b0010100101000010: out_v[162] = 10'b0101001110;
    16'b0010100101000000: out_v[162] = 10'b1101011110;
    16'b0010100101010011: out_v[162] = 10'b1010010000;
    16'b0010100101000001: out_v[162] = 10'b0010011111;
    16'b0000000001010010: out_v[162] = 10'b1100011011;
    16'b0000000001110010: out_v[162] = 10'b0010011100;
    16'b0000000100000001: out_v[162] = 10'b0001011101;
    16'b0010000001110010: out_v[162] = 10'b1010101011;
    16'b0010100100000001: out_v[162] = 10'b1011011110;
    16'b0000000101000010: out_v[162] = 10'b1010110010;
    16'b0000100001000010: out_v[162] = 10'b1011110010;
    16'b0001000101000010: out_v[162] = 10'b1001011000;
    16'b0001000001000010: out_v[162] = 10'b1110101111;
    16'b0001000001000011: out_v[162] = 10'b1010111111;
    16'b0001000001000000: out_v[162] = 10'b0101100010;
    16'b0000100100000000: out_v[162] = 10'b0001111010;
    16'b0000100101000010: out_v[162] = 10'b1001111110;
    16'b0010000101000010: out_v[162] = 10'b1110110000;
    16'b0001100100000000: out_v[162] = 10'b0011110111;
    16'b0010100100000000: out_v[162] = 10'b1010110001;
    16'b0001000001000001: out_v[162] = 10'b0111110011;
    16'b0001100101000010: out_v[162] = 10'b1001001001;
    16'b0000000100000010: out_v[162] = 10'b0110001010;
    16'b0000000100000011: out_v[162] = 10'b1100010110;
    16'b0000100001000001: out_v[162] = 10'b0101101011;
    16'b0001000100000010: out_v[162] = 10'b1101010110;
    16'b0011100101000000: out_v[162] = 10'b0011111000;
    16'b0001000101000000: out_v[162] = 10'b1101101100;
    16'b0011000001000000: out_v[162] = 10'b1111110010;
    16'b0001100101000000: out_v[162] = 10'b0101000111;
    16'b0001000101000001: out_v[162] = 10'b1011100010;
    16'b0011000101000000: out_v[162] = 10'b1110001101;
    16'b0011000101000001: out_v[162] = 10'b1011111011;
    16'b1000000001000010: out_v[162] = 10'b1010101010;
    16'b1000000001000011: out_v[162] = 10'b1111100101;
    default: out_v[162] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001000100000000: out_v[163] = 10'b1010100010;
    16'b0011000000100000: out_v[163] = 10'b1101010111;
    16'b0001000000100000: out_v[163] = 10'b0110101001;
    16'b0000000000101000: out_v[163] = 10'b0001000011;
    16'b0001000000000000: out_v[163] = 10'b0001100111;
    16'b0000000000100000: out_v[163] = 10'b0101001101;
    16'b0010000000100000: out_v[163] = 10'b1111000111;
    16'b0001001000100000: out_v[163] = 10'b1000111010;
    16'b0001000100100000: out_v[163] = 10'b1100111011;
    16'b0001000000101000: out_v[163] = 10'b0000101101;
    16'b0010000000001000: out_v[163] = 10'b0001011111;
    16'b0000000100100000: out_v[163] = 10'b1101010001;
    16'b0010000000101000: out_v[163] = 10'b1010110000;
    16'b0001001000110000: out_v[163] = 10'b1000001011;
    16'b0000000000001000: out_v[163] = 10'b0100001101;
    16'b0000000000000000: out_v[163] = 10'b1010011010;
    16'b0011000000101000: out_v[163] = 10'b0111101110;
    16'b0011000000000000: out_v[163] = 10'b1110000101;
    16'b0010000000000000: out_v[163] = 10'b0000100010;
    16'b0000000100000000: out_v[163] = 10'b0100010010;
    16'b0000001000010000: out_v[163] = 10'b0101010100;
    16'b0001001000010000: out_v[163] = 10'b1001010110;
    16'b0000001100010000: out_v[163] = 10'b0000101111;
    16'b0001000000110000: out_v[163] = 10'b1000110110;
    16'b0001001000000000: out_v[163] = 10'b1001111100;
    16'b0001001000111000: out_v[163] = 10'b1111101110;
    16'b0001010000100000: out_v[163] = 10'b0001100000;
    16'b0011010000101000: out_v[163] = 10'b1100011001;
    16'b0000001000000000: out_v[163] = 10'b1110000011;
    16'b0000001000110000: out_v[163] = 10'b0111110111;
    16'b0001000000100100: out_v[163] = 10'b1101110111;
    16'b0011010000100000: out_v[163] = 10'b1010100111;
    16'b0000001100000000: out_v[163] = 10'b1010001110;
    16'b0100000100000000: out_v[163] = 10'b1010100100;
    16'b0010000100000000: out_v[163] = 10'b0100011011;
    16'b0001010000000000: out_v[163] = 10'b1111100010;
    16'b0000010000000000: out_v[163] = 10'b0010110010;
    16'b0000010000100000: out_v[163] = 10'b0011100100;
    16'b1000000000000000: out_v[163] = 10'b1110000001;
    16'b0100000000000000: out_v[163] = 10'b1011000100;
    16'b0101000100000000: out_v[163] = 10'b0111101011;
    16'b1100000100000000: out_v[163] = 10'b1111011101;
    16'b0011000100000000: out_v[163] = 10'b1101000011;
    16'b0001001100010000: out_v[163] = 10'b0111010101;
    16'b0101000100100000: out_v[163] = 10'b1110000010;
    default: out_v[163] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000000000000: out_v[164] = 10'b1100110000;
    16'b0000100100110000: out_v[164] = 10'b0001100111;
    16'b0000100100110010: out_v[164] = 10'b0011000111;
    16'b0000110101110010: out_v[164] = 10'b1100111011;
    16'b0000100100000000: out_v[164] = 10'b1100110000;
    16'b0000000101000010: out_v[164] = 10'b0011001001;
    16'b0000000100000010: out_v[164] = 10'b0010110011;
    16'b0000000100000000: out_v[164] = 10'b0101011011;
    16'b0000110100110000: out_v[164] = 10'b0100100111;
    16'b0000100100010010: out_v[164] = 10'b1010100101;
    16'b0000100100010000: out_v[164] = 10'b0010111000;
    16'b0000100101110010: out_v[164] = 10'b1000100000;
    16'b0000100000110000: out_v[164] = 10'b1110000110;
    16'b0000000001000000: out_v[164] = 10'b1110011110;
    16'b0000000000010000: out_v[164] = 10'b0110101000;
    16'b0000000100110010: out_v[164] = 10'b0011001111;
    16'b0000000101010010: out_v[164] = 10'b0111001000;
    16'b0000100101010010: out_v[164] = 10'b1010110100;
    16'b0000000101110010: out_v[164] = 10'b1010011100;
    16'b0000000100110000: out_v[164] = 10'b0111010010;
    16'b0000000001000010: out_v[164] = 10'b1111100001;
    16'b0000100001110010: out_v[164] = 10'b0001000001;
    16'b0000110100110010: out_v[164] = 10'b0011000101;
    16'b0000000001110010: out_v[164] = 10'b0101000001;
    16'b0000100000000000: out_v[164] = 10'b1111000011;
    16'b0000000100010000: out_v[164] = 10'b1001100000;
    16'b0000110100010000: out_v[164] = 10'b1011011001;
    16'b0000000001010010: out_v[164] = 10'b1111010011;
    16'b0000100001010010: out_v[164] = 10'b1001001101;
    16'b0000110101010010: out_v[164] = 10'b1001101011;
    16'b0000000100010010: out_v[164] = 10'b0000001101;
    16'b0000110001110010: out_v[164] = 10'b1011111100;
    16'b0000000101000000: out_v[164] = 10'b0001000111;
    16'b0000100101000010: out_v[164] = 10'b0100010111;
    16'b0000110100000000: out_v[164] = 10'b0101000000;
    16'b0000110000110000: out_v[164] = 10'b0101001111;
    16'b0000110000000000: out_v[164] = 10'b0101111010;
    16'b0000110000100000: out_v[164] = 10'b1000100110;
    16'b0000000100000001: out_v[164] = 10'b0001001110;
    16'b0000000100110001: out_v[164] = 10'b0100101101;
    16'b0000000101010000: out_v[164] = 10'b0010111111;
    16'b0000100000010000: out_v[164] = 10'b0000111001;
    16'b0000000101110000: out_v[164] = 10'b0100110010;
    16'b0000000000110000: out_v[164] = 10'b0111111011;
    16'b0000000101110001: out_v[164] = 10'b0001110101;
    16'b0000000000000001: out_v[164] = 10'b1000011100;
    16'b0000110000010000: out_v[164] = 10'b1101100111;
    16'b0000000101000001: out_v[164] = 10'b1010000101;
    16'b0000000001010000: out_v[164] = 10'b1110110010;
    16'b0000000101010001: out_v[164] = 10'b0000010111;
    16'b0000100001110000: out_v[164] = 10'b0110111011;
    16'b0000000001110000: out_v[164] = 10'b1101011101;
    16'b0000100101110000: out_v[164] = 10'b1011001110;
    16'b0000110101110000: out_v[164] = 10'b1011001100;
    16'b0000000000000010: out_v[164] = 10'b1011010101;
    16'b0000000100010001: out_v[164] = 10'b1110010110;
    16'b0000100100110001: out_v[164] = 10'b0100110111;
    16'b0000110001110000: out_v[164] = 10'b0100110110;
    16'b0000100001010000: out_v[164] = 10'b1010100100;
    16'b0000110100100000: out_v[164] = 10'b0101101111;
    16'b0000000000100000: out_v[164] = 10'b1001001101;
    16'b0000100100100000: out_v[164] = 10'b0010011000;
    16'b0000000100100000: out_v[164] = 10'b1100100100;
    16'b0000000000110001: out_v[164] = 10'b1101110111;
    16'b0000000001110001: out_v[164] = 10'b1001001110;
    16'b0000000001000001: out_v[164] = 10'b0110101010;
    16'b0000100000000010: out_v[164] = 10'b0001110111;
    16'b0000110000000010: out_v[164] = 10'b1010110010;
    16'b0000100001000000: out_v[164] = 10'b0101111011;
    16'b0000100100000010: out_v[164] = 10'b1110111101;
    16'b0000110100000010: out_v[164] = 10'b1000100011;
    16'b0000110001000000: out_v[164] = 10'b1111100000;
    16'b0000010100000000: out_v[164] = 10'b0101001001;
    16'b0000000101000011: out_v[164] = 10'b1011100010;
    16'b0000100000100000: out_v[164] = 10'b1011001110;
    default: out_v[164] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1000010000000000: out_v[165] = 10'b0011000011;
    16'b1001110000000000: out_v[165] = 10'b0001000111;
    16'b1001010000000000: out_v[165] = 10'b0001110101;
    16'b0000010000000000: out_v[165] = 10'b1111010011;
    16'b0001100000000000: out_v[165] = 10'b0110110101;
    16'b1001010100000000: out_v[165] = 10'b0100111100;
    16'b1001000000000000: out_v[165] = 10'b0100110001;
    16'b0001010000000000: out_v[165] = 10'b0001001111;
    16'b0001110000000000: out_v[165] = 10'b1010010111;
    16'b1001010000000001: out_v[165] = 10'b1000000110;
    16'b1001010001000000: out_v[165] = 10'b1101011000;
    16'b0001000001000000: out_v[165] = 10'b0100010011;
    16'b0001000000000000: out_v[165] = 10'b0101110101;
    16'b1001110000000001: out_v[165] = 10'b1101000110;
    16'b1001000001000000: out_v[165] = 10'b0111111010;
    16'b1001110100000000: out_v[165] = 10'b0100101000;
    16'b0000000000000000: out_v[165] = 10'b1010001001;
    16'b1000110000000001: out_v[165] = 10'b1110011101;
    16'b0001000010000000: out_v[165] = 10'b1010101111;
    16'b1000000000000000: out_v[165] = 10'b1001100111;
    16'b1001100000000000: out_v[165] = 10'b1001110111;
    16'b1001110001000000: out_v[165] = 10'b1111101011;
    16'b1000010100000000: out_v[165] = 10'b1000011001;
    16'b1001000100000000: out_v[165] = 10'b1110110011;
    16'b0001000100000000: out_v[165] = 10'b0110001110;
    16'b0000000100000000: out_v[165] = 10'b0000010110;
    16'b1000000100000000: out_v[165] = 10'b1001010100;
    16'b0001000100000001: out_v[165] = 10'b0111010110;
    16'b0000000110000000: out_v[165] = 10'b1001110110;
    16'b0001000110000000: out_v[165] = 10'b0100000110;
    16'b0001010100000000: out_v[165] = 10'b1011011110;
    16'b0000010010000000: out_v[165] = 10'b0001110110;
    16'b0001010110000000: out_v[165] = 10'b0000100101;
    16'b0001010010000000: out_v[165] = 10'b1000100101;
    16'b0000010100000000: out_v[165] = 10'b1110100111;
    16'b0000000010000000: out_v[165] = 10'b0101010001;
    16'b0000010110000000: out_v[165] = 10'b1111010010;
    16'b1001010110000000: out_v[165] = 10'b0010001011;
    16'b1000010110000000: out_v[165] = 10'b1110000011;
    16'b1001100000000001: out_v[165] = 10'b0110101110;
    16'b0001010100000001: out_v[165] = 10'b0110011110;
    16'b1000010010000000: out_v[165] = 10'b1101011100;
    16'b0000010100000001: out_v[165] = 10'b1101011101;
    16'b0001110100000000: out_v[165] = 10'b1010011001;
    16'b1001000100000001: out_v[165] = 10'b1011010010;
    16'b1001000110000000: out_v[165] = 10'b1010001110;
    16'b0000010110000001: out_v[165] = 10'b1011001000;
    16'b1000010100000001: out_v[165] = 10'b1001000010;
    16'b0000000100000001: out_v[165] = 10'b0000011010;
    16'b1000000110000000: out_v[165] = 10'b0010011001;
    16'b1001010100000001: out_v[165] = 10'b0101110100;
    16'b0001010110000001: out_v[165] = 10'b1111110111;
    16'b1000110100000000: out_v[165] = 10'b0011101010;
    16'b1000100000000000: out_v[165] = 10'b0010101010;
    16'b0000100000000000: out_v[165] = 10'b0000110111;
    16'b1000100100000000: out_v[165] = 10'b1100000111;
    16'b0000100100000000: out_v[165] = 10'b1100110111;
    16'b1000110000000000: out_v[165] = 10'b0011110011;
    16'b0000010011000000: out_v[165] = 10'b0000010111;
    16'b0000010101000000: out_v[165] = 10'b0111010111;
    16'b0000110000000000: out_v[165] = 10'b1110010110;
    16'b0000010111000000: out_v[165] = 10'b0101110001;
    16'b0000010001000000: out_v[165] = 10'b1100111010;
    16'b1011100000000000: out_v[165] = 10'b1100101110;
    16'b1001100100000000: out_v[165] = 10'b1100010100;
    16'b0001100100000000: out_v[165] = 10'b1001110011;
    16'b0100010110000000: out_v[165] = 10'b0011111011;
    16'b0000000000000100: out_v[165] = 10'b1111110100;
    16'b0000010000000100: out_v[165] = 10'b0101001010;
    16'b1000010100000100: out_v[165] = 10'b1101011010;
    16'b1000010000000100: out_v[165] = 10'b1010111011;
    16'b0000000100000100: out_v[165] = 10'b1100001111;
    16'b0000010100000100: out_v[165] = 10'b0010101111;
    16'b1000010001000000: out_v[165] = 10'b0100010011;
    16'b1000000010000000: out_v[165] = 10'b0100101001;
    16'b1000010101000000: out_v[165] = 10'b1010000111;
    16'b1000000001000000: out_v[165] = 10'b1100001100;
    16'b1000000101000000: out_v[165] = 10'b0001110100;
    16'b1001100100000001: out_v[165] = 10'b0010111100;
    default: out_v[165] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010011001110000: out_v[166] = 10'b0101110111;
    16'b0010000000000000: out_v[166] = 10'b0111001101;
    16'b0010000000010000: out_v[166] = 10'b1100011011;
    16'b0010010000010000: out_v[166] = 10'b1001000101;
    16'b0010011000010000: out_v[166] = 10'b1001000100;
    16'b0010000000000100: out_v[166] = 10'b0011011000;
    16'b0010000001000000: out_v[166] = 10'b1010111100;
    16'b0000000000000100: out_v[166] = 10'b0011100011;
    16'b0010010000000100: out_v[166] = 10'b0011000111;
    16'b0010001001000100: out_v[166] = 10'b1111000011;
    16'b0010011000110000: out_v[166] = 10'b1110100000;
    16'b0010011001000000: out_v[166] = 10'b0100000010;
    16'b0010010000010100: out_v[166] = 10'b0001000001;
    16'b0010010000000000: out_v[166] = 10'b0001010111;
    16'b0010011001000100: out_v[166] = 10'b1011000010;
    16'b0010000000010100: out_v[166] = 10'b0111101001;
    16'b0010011001010100: out_v[166] = 10'b0001100000;
    16'b0000010100110000: out_v[166] = 10'b0010111110;
    16'b0010000001000100: out_v[166] = 10'b1000111101;
    16'b0010001000000100: out_v[166] = 10'b0111011111;
    16'b0000000000000000: out_v[166] = 10'b0111001101;
    16'b0010011000010100: out_v[166] = 10'b0001101111;
    16'b0010010100110000: out_v[166] = 10'b0000101011;
    16'b0000010000010000: out_v[166] = 10'b0011001011;
    16'b0000001001000000: out_v[166] = 10'b0001000111;
    16'b0010010000110000: out_v[166] = 10'b0111100011;
    16'b0010011000000100: out_v[166] = 10'b1111011010;
    16'b0000011001000000: out_v[166] = 10'b0111010001;
    16'b0010001001000000: out_v[166] = 10'b0011010011;
    16'b0000001001000100: out_v[166] = 10'b0001100011;
    16'b0000011000010100: out_v[166] = 10'b0001010101;
    16'b0000010000010100: out_v[166] = 10'b1011100010;
    16'b0010011001010000: out_v[166] = 10'b0100110110;
    16'b0010011000000000: out_v[166] = 10'b0001011110;
    16'b0000010000110000: out_v[166] = 10'b1000101001;
    16'b0000010000000000: out_v[166] = 10'b1100011001;
    16'b0000001000000100: out_v[166] = 10'b1100100110;
    16'b0000010000100000: out_v[166] = 10'b0010011110;
    16'b0000001000000000: out_v[166] = 10'b1100000110;
    16'b0000010000000100: out_v[166] = 10'b0010000011;
    16'b0000000000100000: out_v[166] = 10'b0010100010;
    16'b0000101000000000: out_v[166] = 10'b1110111111;
    16'b0000000000100100: out_v[166] = 10'b0011101011;
    16'b0000000000010000: out_v[166] = 10'b0111110011;
    16'b0000010000100100: out_v[166] = 10'b0101010000;
    16'b0010010001010100: out_v[166] = 10'b1010101000;
    16'b0000011000000100: out_v[166] = 10'b0111001000;
    16'b0000010001010100: out_v[166] = 10'b0010101010;
    16'b0000010100010100: out_v[166] = 10'b1001111100;
    16'b0000011001010100: out_v[166] = 10'b1000010101;
    16'b0000000000010100: out_v[166] = 10'b0110110101;
    16'b0000011001000100: out_v[166] = 10'b0001000111;
    16'b0000011001010110: out_v[166] = 10'b0010111110;
    16'b0000011000000000: out_v[166] = 10'b1011101100;
    16'b0000011000010000: out_v[166] = 10'b1111000101;
    16'b0000011000000110: out_v[166] = 10'b1111111010;
    16'b0000011000010010: out_v[166] = 10'b1110110111;
    16'b0000000001000100: out_v[166] = 10'b1101010100;
    16'b0000000001000000: out_v[166] = 10'b1000111100;
    16'b0000011000010110: out_v[166] = 10'b1010001001;
    16'b0000001000010100: out_v[166] = 10'b1111111000;
    16'b0010001000000000: out_v[166] = 10'b1101011110;
    16'b0000010001000100: out_v[166] = 10'b0100111101;
    16'b0010001000010000: out_v[166] = 10'b0101010100;
    16'b0000011001010000: out_v[166] = 10'b0101000110;
    16'b0010010001000100: out_v[166] = 10'b0100110111;
    16'b0000011100010100: out_v[166] = 10'b1011000110;
    16'b0000010000010110: out_v[166] = 10'b0000011110;
    16'b0010010001110000: out_v[166] = 10'b1011010110;
    16'b0000010001000000: out_v[166] = 10'b0010111000;
    16'b0000011001110000: out_v[166] = 10'b1010010100;
    16'b0000010101110000: out_v[166] = 10'b1111010000;
    16'b0010010001000000: out_v[166] = 10'b0101100100;
    16'b0000010001010000: out_v[166] = 10'b1001011100;
    16'b0000010001100000: out_v[166] = 10'b0000001001;
    16'b0010010101110000: out_v[166] = 10'b0010011101;
    16'b0000010001110000: out_v[166] = 10'b1011001100;
    16'b0010010001010000: out_v[166] = 10'b1011000101;
    16'b0000001100000000: out_v[166] = 10'b0001111010;
    16'b0000000001010000: out_v[166] = 10'b0011111101;
    16'b0000000101000000: out_v[166] = 10'b0001110111;
    16'b0000000101010000: out_v[166] = 10'b1101011111;
    16'b0010001100000000: out_v[166] = 10'b1110110000;
    16'b0000001000110000: out_v[166] = 10'b0011110000;
    16'b0000000001100000: out_v[166] = 10'b1001011101;
    16'b0000000001010100: out_v[166] = 10'b0010110010;
    16'b0010001001010000: out_v[166] = 10'b1101000111;
    16'b0010001000110000: out_v[166] = 10'b0111010010;
    16'b0000001000010000: out_v[166] = 10'b0111111010;
    16'b0000100001000100: out_v[166] = 10'b1010100011;
    16'b0010001101000000: out_v[166] = 10'b0101111001;
    16'b0000000100000000: out_v[166] = 10'b0111110001;
    16'b0010000101000000: out_v[166] = 10'b0001111111;
    16'b0000001001100000: out_v[166] = 10'b1111000000;
    16'b0000000000110000: out_v[166] = 10'b0100011110;
    16'b0000101000000100: out_v[166] = 10'b0010111000;
    16'b0000001100010000: out_v[166] = 10'b0000011001;
    16'b0000011000110000: out_v[166] = 10'b1001100011;
    16'b0000000001110000: out_v[166] = 10'b0000110110;
    16'b0000001101000000: out_v[166] = 10'b0110001101;
    16'b0010001100010000: out_v[166] = 10'b1101100010;
    16'b0010000001110000: out_v[166] = 10'b1001100100;
    16'b0000001001110000: out_v[166] = 10'b0110010111;
    16'b0010000001100000: out_v[166] = 10'b1101010011;
    16'b0000001000100000: out_v[166] = 10'b1101000100;
    16'b0010000001010000: out_v[166] = 10'b1100011101;
    16'b0010001000100000: out_v[166] = 10'b0110010010;
    16'b0000100000000000: out_v[166] = 10'b0011110011;
    16'b0000100000000100: out_v[166] = 10'b1100101000;
    16'b0000100001000000: out_v[166] = 10'b1111010000;
    16'b0010001001010100: out_v[166] = 10'b0010011111;
    16'b0010001000010100: out_v[166] = 10'b0011101111;
    16'b0010000000100000: out_v[166] = 10'b0110001110;
    16'b0010000100000000: out_v[166] = 10'b0111100000;
    16'b0000000010000000: out_v[166] = 10'b1010001111;
    16'b0000010000110100: out_v[166] = 10'b0111000111;
    16'b0010000000110000: out_v[166] = 10'b0111110010;
    16'b0000000000110100: out_v[166] = 10'b0010010101;
    16'b0000000100100000: out_v[166] = 10'b0010101111;
    16'b0010000100100000: out_v[166] = 10'b0011010111;
    16'b0000000100110000: out_v[166] = 10'b0111011001;
    16'b0000011001100000: out_v[166] = 10'b0110110010;
    16'b0000010101110100: out_v[166] = 10'b0011111000;
    16'b0000011000100000: out_v[166] = 10'b1101110111;
    16'b0010011101110000: out_v[166] = 10'b0110000010;
    16'b0000011000110100: out_v[166] = 10'b1100111110;
    16'b0000101001000000: out_v[166] = 10'b1001011010;
    16'b0000011100110000: out_v[166] = 10'b1110101010;
    16'b0000011101110000: out_v[166] = 10'b1111011011;
    16'b0000010100110100: out_v[166] = 10'b0101110111;
    16'b0000010001110100: out_v[166] = 10'b0101000001;
    16'b0000011101110100: out_v[166] = 10'b1000011110;
    16'b0000011001110100: out_v[166] = 10'b1110100110;
    16'b0000000001100100: out_v[166] = 10'b0100001001;
    16'b0000011100010000: out_v[166] = 10'b1011100110;
    16'b0010011100010000: out_v[166] = 10'b1000100100;
    16'b0000010101010000: out_v[166] = 10'b1111001101;
    16'b0000010100010000: out_v[166] = 10'b1011000011;
    default: out_v[166] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000000010000: out_v[167] = 10'b0010110011;
    16'b0000000000010010: out_v[167] = 10'b0101011011;
    16'b0010000000010010: out_v[167] = 10'b0000011001;
    16'b0010000000000010: out_v[167] = 10'b1000001011;
    16'b0010000000110010: out_v[167] = 10'b1011010101;
    16'b0000000000000010: out_v[167] = 10'b0000100111;
    16'b0010000000000000: out_v[167] = 10'b0010110011;
    16'b0000000000110000: out_v[167] = 10'b0010010110;
    16'b0000000000010011: out_v[167] = 10'b0010101101;
    16'b0000000001110011: out_v[167] = 10'b0111101111;
    16'b0000000001010010: out_v[167] = 10'b0000001010;
    16'b0000000000110010: out_v[167] = 10'b1001010011;
    16'b0010010000010010: out_v[167] = 10'b0001001001;
    16'b0000000001110010: out_v[167] = 10'b1000101000;
    16'b0000000000010001: out_v[167] = 10'b1000100001;
    16'b0010000000010000: out_v[167] = 10'b0010100011;
    16'b0010010000000010: out_v[167] = 10'b0110000111;
    16'b0000000001010011: out_v[167] = 10'b0100100101;
    16'b0010000001010010: out_v[167] = 10'b1011110110;
    16'b0000000000110011: out_v[167] = 10'b0000100110;
    16'b0000000000000000: out_v[167] = 10'b0110100011;
    16'b0000000000110001: out_v[167] = 10'b1101010110;
    16'b0000000000000001: out_v[167] = 10'b1000101011;
    16'b0000000001110001: out_v[167] = 10'b1000100010;
    16'b0000000001000000: out_v[167] = 10'b1001001010;
    16'b0000000001000001: out_v[167] = 10'b0110101110;
    16'b0000000001100001: out_v[167] = 10'b0111110100;
    16'b0000000001010001: out_v[167] = 10'b0101110101;
    16'b0000000001100000: out_v[167] = 10'b1110110011;
    16'b0000000001010000: out_v[167] = 10'b1001011101;
    16'b0000000000100000: out_v[167] = 10'b0111001110;
    16'b0000010000110011: out_v[167] = 10'b1101011110;
    16'b0000000000100001: out_v[167] = 10'b1000111101;
    16'b0010010001000001: out_v[167] = 10'b1101010101;
    16'b0000000000100011: out_v[167] = 10'b0100100111;
    16'b0000010000100001: out_v[167] = 10'b0110010011;
    16'b0000000000111011: out_v[167] = 10'b1001001001;
    16'b0000000000100010: out_v[167] = 10'b1111010010;
    16'b0000000001000011: out_v[167] = 10'b1011001100;
    16'b0000000001100011: out_v[167] = 10'b0000011100;
    16'b0000010000100000: out_v[167] = 10'b1100100110;
    16'b0010000001000001: out_v[167] = 10'b1111001110;
    16'b0010000000110000: out_v[167] = 10'b0011011010;
    16'b0010000000110011: out_v[167] = 10'b0110001111;
    16'b0010000000100011: out_v[167] = 10'b0100110100;
    16'b0010010000110010: out_v[167] = 10'b0011101010;
    16'b0010000000100010: out_v[167] = 10'b0101001100;
    16'b0010000001010011: out_v[167] = 10'b1110011110;
    16'b0000010000110010: out_v[167] = 10'b0111001000;
    16'b0000000000111010: out_v[167] = 10'b1111110111;
    16'b0010010001100001: out_v[167] = 10'b0010011110;
    16'b0000010001000001: out_v[167] = 10'b1001000110;
    16'b0010000001100001: out_v[167] = 10'b0111001101;
    16'b0010000000100001: out_v[167] = 10'b1100111010;
    16'b0010000000100000: out_v[167] = 10'b0111000010;
    16'b0000000001011010: out_v[167] = 10'b1101001001;
    16'b0000000001011000: out_v[167] = 10'b1111110011;
    16'b0000010001100001: out_v[167] = 10'b1010101010;
    16'b0000000001110000: out_v[167] = 10'b1100110000;
    16'b0000010001000000: out_v[167] = 10'b1100011011;
    16'b0000010001110001: out_v[167] = 10'b0101011011;
    16'b0000000001000010: out_v[167] = 10'b1010101011;
    16'b0000000001111011: out_v[167] = 10'b1010000101;
    16'b0000000001111010: out_v[167] = 10'b0111011011;
    16'b0010010001110001: out_v[167] = 10'b0100010010;
    16'b0000010001010010: out_v[167] = 10'b0111011011;
    16'b0000010001010001: out_v[167] = 10'b1100110011;
    16'b0000010001000010: out_v[167] = 10'b0111001010;
    16'b0000000001111001: out_v[167] = 10'b1111000011;
    16'b0010000001010001: out_v[167] = 10'b0111010001;
    16'b0000010001010011: out_v[167] = 10'b1000011011;
    16'b0010000001110001: out_v[167] = 10'b0110011001;
    16'b0000000001100010: out_v[167] = 10'b1010100010;
    16'b0000000011000000: out_v[167] = 10'b1011001010;
    16'b0000000001011011: out_v[167] = 10'b0110110010;
    16'b0010000001110011: out_v[167] = 10'b0101011101;
    16'b0010000000110001: out_v[167] = 10'b1101010000;
    16'b0010010000100001: out_v[167] = 10'b0110011011;
    16'b0010000000000001: out_v[167] = 10'b1100100011;
    16'b0010000001100000: out_v[167] = 10'b1000011011;
    16'b0010010000110001: out_v[167] = 10'b1110100000;
    16'b0000010000110001: out_v[167] = 10'b0111111011;
    16'b0010000001110000: out_v[167] = 10'b1001110110;
    16'b0010000001010000: out_v[167] = 10'b1101110000;
    16'b0010000001110010: out_v[167] = 10'b0011110101;
    16'b0010010001000000: out_v[167] = 10'b1000100010;
    16'b0010000000010001: out_v[167] = 10'b1001100110;
    16'b0010000001000000: out_v[167] = 10'b1010111101;
    16'b0010000001000010: out_v[167] = 10'b1110100101;
    16'b0010010001010010: out_v[167] = 10'b0010100000;
    16'b0000000000000011: out_v[167] = 10'b0111010011;
    16'b0010000000000011: out_v[167] = 10'b0101111010;
    16'b0010000001000011: out_v[167] = 10'b0111011010;
    16'b0010010000110000: out_v[167] = 10'b1001000110;
    16'b0010010001100000: out_v[167] = 10'b0110001011;
    16'b0010010001110000: out_v[167] = 10'b1111000011;
    16'b0010010000100000: out_v[167] = 10'b0100011000;
    16'b0010010000000000: out_v[167] = 10'b0110010111;
    16'b0000010000110000: out_v[167] = 10'b1010100111;
    16'b0000010000000000: out_v[167] = 10'b1011110101;
    16'b0010000000010011: out_v[167] = 10'b1010000111;
    default: out_v[167] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010001100000000: out_v[168] = 10'b0000000101;
    16'b0010011001011000: out_v[168] = 10'b1011100111;
    16'b0010001101011001: out_v[168] = 10'b0010011001;
    16'b0000001101000000: out_v[168] = 10'b0110000111;
    16'b0010001000000000: out_v[168] = 10'b0110000101;
    16'b0010001001011000: out_v[168] = 10'b0001101000;
    16'b0000001001011000: out_v[168] = 10'b1001000011;
    16'b0000000001010001: out_v[168] = 10'b1100011101;
    16'b0000001101011000: out_v[168] = 10'b0110101111;
    16'b0000011001011001: out_v[168] = 10'b1111101110;
    16'b0000000101011000: out_v[168] = 10'b0101011011;
    16'b0000000001010000: out_v[168] = 10'b1000001111;
    16'b0010000000000000: out_v[168] = 10'b1010001010;
    16'b0010000101000000: out_v[168] = 10'b0100111010;
    16'b0000000101011001: out_v[168] = 10'b1110010110;
    16'b0010001001000000: out_v[168] = 10'b0011001100;
    16'b0000010101011000: out_v[168] = 10'b1110011110;
    16'b0010001101011000: out_v[168] = 10'b0011000001;
    16'b0010000001000000: out_v[168] = 10'b0010001111;
    16'b0000011101011000: out_v[168] = 10'b1011011100;
    16'b0010000101011000: out_v[168] = 10'b1110100110;
    16'b0010001001000001: out_v[168] = 10'b0100001101;
    16'b0000000001000000: out_v[168] = 10'b1110010111;
    16'b0010001101000000: out_v[168] = 10'b0101000111;
    16'b0010001101001000: out_v[168] = 10'b1110001011;
    16'b0000000001011000: out_v[168] = 10'b1010010011;
    16'b0000000101010000: out_v[168] = 10'b1100000111;
    16'b0000001101011001: out_v[168] = 10'b0110011101;
    16'b0000001001010001: out_v[168] = 10'b0110110111;
    16'b0000000001011001: out_v[168] = 10'b0001011110;
    16'b0000001001011001: out_v[168] = 10'b0010100011;
    16'b0010001101010000: out_v[168] = 10'b0011101110;
    16'b0000001001010000: out_v[168] = 10'b0111001101;
    16'b0010000001011000: out_v[168] = 10'b1011100001;
    16'b0000001001000001: out_v[168] = 10'b1110011101;
    16'b0010001001010001: out_v[168] = 10'b1001111010;
    16'b0000011101011001: out_v[168] = 10'b1001110101;
    16'b0010001100001000: out_v[168] = 10'b0100000101;
    16'b0000001101010000: out_v[168] = 10'b1010011111;
    16'b0000000101000000: out_v[168] = 10'b0100010011;
    16'b0000001101010001: out_v[168] = 10'b0000010111;
    16'b0010000100000000: out_v[168] = 10'b1110010100;
    16'b0000011001011000: out_v[168] = 10'b0101011110;
    16'b0010001001010000: out_v[168] = 10'b1011100010;
    16'b0000000001000001: out_v[168] = 10'b0110010101;
    16'b0010001001011001: out_v[168] = 10'b1001110101;
    16'b0010000101010000: out_v[168] = 10'b0111101010;
    16'b0010001000000001: out_v[168] = 10'b1000000010;
    16'b0000000000000000: out_v[168] = 10'b0110110110;
    16'b0000000100000000: out_v[168] = 10'b0010011010;
    16'b0000001000000000: out_v[168] = 10'b0001010010;
    16'b0000001100000000: out_v[168] = 10'b1000111100;
    16'b0010000000000001: out_v[168] = 10'b0100001001;
    16'b0000001000000001: out_v[168] = 10'b1001000000;
    16'b0010000100000001: out_v[168] = 10'b1100000011;
    16'b0000001101000001: out_v[168] = 10'b1110000110;
    16'b0010001101000001: out_v[168] = 10'b1011011100;
    16'b0010001100000001: out_v[168] = 10'b1010011111;
    16'b0000000100001000: out_v[168] = 10'b0101101000;
    16'b0010000101000001: out_v[168] = 10'b0100001001;
    16'b0010000100001000: out_v[168] = 10'b1001000111;
    16'b0010001100010000: out_v[168] = 10'b1000011110;
    16'b0000000100000001: out_v[168] = 10'b1011110110;
    16'b0010000000001000: out_v[168] = 10'b1010011010;
    16'b0000000000001000: out_v[168] = 10'b1000110111;
    16'b0010000001001000: out_v[168] = 10'b0000010101;
    16'b0010001000001001: out_v[168] = 10'b0100110010;
    16'b0010000101001000: out_v[168] = 10'b1110001011;
    16'b0010001001001000: out_v[168] = 10'b0110001101;
    16'b0010000000001001: out_v[168] = 10'b1011110010;
    16'b0010000000010000: out_v[168] = 10'b0011010010;
    16'b0000000001001000: out_v[168] = 10'b1011010111;
    16'b0010000001001001: out_v[168] = 10'b1001110010;
    16'b0010000000011000: out_v[168] = 10'b0111111110;
    16'b1010001011001000: out_v[168] = 10'b0011101010;
    16'b0010001000001000: out_v[168] = 10'b1110111100;
    16'b0010000000011001: out_v[168] = 10'b1011100110;
    16'b0000000000010000: out_v[168] = 10'b0010100110;
    16'b0010100000001000: out_v[168] = 10'b1001000111;
    16'b0010011001000000: out_v[168] = 10'b0000100100;
    16'b0000000000000001: out_v[168] = 10'b0011100100;
    16'b1000001010000000: out_v[168] = 10'b1000110110;
    16'b0000001100000001: out_v[168] = 10'b1010110010;
    16'b0000000010000001: out_v[168] = 10'b0011001110;
    16'b0000001000001000: out_v[168] = 10'b1100110110;
    16'b1000001000000000: out_v[168] = 10'b0000111100;
    16'b0000010000000000: out_v[168] = 10'b0100101101;
    16'b1000000010000001: out_v[168] = 10'b1011111010;
    16'b1000001010000001: out_v[168] = 10'b0000111101;
    16'b0010010001000000: out_v[168] = 10'b0111100000;
    16'b0000000100001001: out_v[168] = 10'b0001100100;
    16'b1000000010000000: out_v[168] = 10'b1011111010;
    16'b0000011000000000: out_v[168] = 10'b1001111010;
    16'b0000001100001000: out_v[168] = 10'b0001100010;
    16'b1000000000001000: out_v[168] = 10'b0000010110;
    16'b1000000000000000: out_v[168] = 10'b0010111111;
    16'b0000000000001001: out_v[168] = 10'b0110101000;
    16'b0010011000000000: out_v[168] = 10'b1001110010;
    16'b0000001100001001: out_v[168] = 10'b0001011110;
    16'b0010001100011000: out_v[168] = 10'b0011001110;
    16'b0000001100010000: out_v[168] = 10'b1110000110;
    16'b0000001100011000: out_v[168] = 10'b1111000000;
    16'b0000001000011000: out_v[168] = 10'b1000110100;
    16'b0010001000010000: out_v[168] = 10'b0111110110;
    16'b0000001000010000: out_v[168] = 10'b0100111011;
    16'b0000001000001001: out_v[168] = 10'b1011100000;
    16'b0010000001010000: out_v[168] = 10'b1111000110;
    16'b0000001001000000: out_v[168] = 10'b1110000110;
    16'b0010011101000000: out_v[168] = 10'b1100110101;
    16'b0010000001000001: out_v[168] = 10'b0100011010;
    16'b0010010101000000: out_v[168] = 10'b1010111110;
    default: out_v[168] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000000001100: out_v[169] = 10'b1110100010;
    16'b1000000001001000: out_v[169] = 10'b1010110100;
    16'b1000000001001010: out_v[169] = 10'b0000011111;
    16'b0000000000001010: out_v[169] = 10'b1100101011;
    16'b0000000000000000: out_v[169] = 10'b0001111101;
    16'b0000000000000010: out_v[169] = 10'b1100000011;
    16'b0000000000001000: out_v[169] = 10'b1001001111;
    16'b0000000001001010: out_v[169] = 10'b0000001011;
    16'b0000000001001000: out_v[169] = 10'b1000011011;
    16'b0000000001001110: out_v[169] = 10'b1000010101;
    16'b0000000000001110: out_v[169] = 10'b1010110110;
    16'b0000000001000010: out_v[169] = 10'b0101001111;
    16'b1000000001001110: out_v[169] = 10'b1011100100;
    16'b1000000001000000: out_v[169] = 10'b1000011101;
    16'b0000000000000110: out_v[169] = 10'b0010100001;
    16'b0000000001000110: out_v[169] = 10'b0000000111;
    16'b0000000001000000: out_v[169] = 10'b1100100001;
    16'b1000000001000010: out_v[169] = 10'b1000110011;
    16'b0000000001001100: out_v[169] = 10'b1100100110;
    16'b1100000001000000: out_v[169] = 10'b1010100011;
    16'b0000000010000000: out_v[169] = 10'b0110110010;
    16'b0000000011000000: out_v[169] = 10'b1100100100;
    16'b0000000010001100: out_v[169] = 10'b0100010010;
    16'b1000000011000000: out_v[169] = 10'b1111000000;
    16'b0000000010000100: out_v[169] = 10'b1001000110;
    16'b0000000010001000: out_v[169] = 10'b1001100100;
    16'b1100000011000000: out_v[169] = 10'b1100011010;
    16'b0000010011000000: out_v[169] = 10'b1011100111;
    16'b0000000011001100: out_v[169] = 10'b0010010010;
    16'b0000000011001000: out_v[169] = 10'b0011011010;
    16'b0000010010000000: out_v[169] = 10'b1111101110;
    16'b0000000010001010: out_v[169] = 10'b1001110111;
    16'b0001000010000000: out_v[169] = 10'b0010100011;
    16'b1000000011001100: out_v[169] = 10'b1010001110;
    16'b1000010011001000: out_v[169] = 10'b0011111011;
    16'b1000000011001000: out_v[169] = 10'b0010011011;
    16'b0000000010000010: out_v[169] = 10'b0001111111;
    16'b1000000001001100: out_v[169] = 10'b0111011110;
    16'b0000000011000010: out_v[169] = 10'b1010011110;
    16'b1000000011001010: out_v[169] = 10'b0011001111;
    16'b0001000010001000: out_v[169] = 10'b1111010111;
    16'b0001001010001100: out_v[169] = 10'b1011101010;
    16'b0001000010001100: out_v[169] = 10'b1011011100;
    16'b0001001010001000: out_v[169] = 10'b1001100101;
    16'b1000000011001110: out_v[169] = 10'b1110110010;
    16'b1000000011000100: out_v[169] = 10'b1100001101;
    16'b0000010010001100: out_v[169] = 10'b1011000010;
    16'b0000000010001110: out_v[169] = 10'b0101110000;
    16'b0000010010001000: out_v[169] = 10'b1111100001;
    16'b0000010011001000: out_v[169] = 10'b1010100111;
    16'b1000000011000010: out_v[169] = 10'b1101001100;
    16'b0001000000000100: out_v[169] = 10'b1001101101;
    16'b0000000110000000: out_v[169] = 10'b1010110000;
    16'b0001000011001100: out_v[169] = 10'b0010101000;
    16'b0000000110001100: out_v[169] = 10'b0100101010;
    16'b1000000010001000: out_v[169] = 10'b1110011011;
    16'b0001000000001100: out_v[169] = 10'b1101000101;
    16'b0001000010000100: out_v[169] = 10'b1000011110;
    16'b1000000010000000: out_v[169] = 10'b0011011000;
    16'b1000000000001100: out_v[169] = 10'b1010011100;
    16'b1001000001001100: out_v[169] = 10'b0100110010;
    16'b1001000011001100: out_v[169] = 10'b1000001001;
    16'b0001000001001100: out_v[169] = 10'b1101000001;
    16'b1000000000001000: out_v[169] = 10'b0101100001;
    16'b0001001000001100: out_v[169] = 10'b0111010010;
    16'b0000000110001000: out_v[169] = 10'b1001110111;
    16'b1000000000000000: out_v[169] = 10'b0011001111;
    16'b1001000010001100: out_v[169] = 10'b0101110111;
    16'b1000000010001100: out_v[169] = 10'b1001101001;
    16'b0000000110000010: out_v[169] = 10'b1010000001;
    16'b0100000010000010: out_v[169] = 10'b0001110110;
    16'b0001000010000010: out_v[169] = 10'b0110111011;
    16'b0100000010000000: out_v[169] = 10'b1111011010;
    16'b0001000010001110: out_v[169] = 10'b0100110110;
    16'b0000000010000110: out_v[169] = 10'b0110000010;
    16'b0100000000000010: out_v[169] = 10'b0100011110;
    16'b0000000011001010: out_v[169] = 10'b0010110101;
    16'b1100000001001010: out_v[169] = 10'b1010001100;
    16'b0000000100000000: out_v[169] = 10'b1011000010;
    16'b0000000100000010: out_v[169] = 10'b1010100010;
    16'b0100000011000000: out_v[169] = 10'b1011001110;
    16'b1100000001001000: out_v[169] = 10'b1010110001;
    16'b0100000010001110: out_v[169] = 10'b0100101101;
    16'b1100000011001110: out_v[169] = 10'b1001110111;
    16'b0000000011001110: out_v[169] = 10'b1011000010;
    16'b0100000001000000: out_v[169] = 10'b1001010100;
    16'b0000000110001110: out_v[169] = 10'b0101011000;
    16'b1100000001001110: out_v[169] = 10'b1011110110;
    16'b0100000011001110: out_v[169] = 10'b1010110110;
    16'b0000000110001010: out_v[169] = 10'b0100111101;
    16'b1100000011001000: out_v[169] = 10'b1101010010;
    16'b0000000010101010: out_v[169] = 10'b0110100001;
    16'b0000000010100000: out_v[169] = 10'b1011000010;
    16'b0000010010001010: out_v[169] = 10'b1111101100;
    16'b0000000010101000: out_v[169] = 10'b1100101101;
    16'b0000010010101010: out_v[169] = 10'b1001101111;
    16'b0000001010001010: out_v[169] = 10'b1111011001;
    16'b0000000000101010: out_v[169] = 10'b1011000100;
    16'b0000000000101000: out_v[169] = 10'b0011001100;
    16'b0000000010100010: out_v[169] = 10'b0111111111;
    16'b0000000000100000: out_v[169] = 10'b0101000010;
    16'b0000010010001110: out_v[169] = 10'b1001111010;
    16'b0000010000001010: out_v[169] = 10'b1111001010;
    16'b0001000000000000: out_v[169] = 10'b0111010011;
    16'b0001000100000000: out_v[169] = 10'b1000110101;
    16'b0000000000001111: out_v[169] = 10'b0110010110;
    16'b0000000100001010: out_v[169] = 10'b1111011110;
    16'b0001000110000000: out_v[169] = 10'b1000110011;
    16'b0000100010001110: out_v[169] = 10'b1011101111;
    default: out_v[169] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001000010000000: out_v[170] = 10'b1100000111;
    16'b0001000111010000: out_v[170] = 10'b0001000011;
    16'b0001000101110010: out_v[170] = 10'b1011011110;
    16'b0001000011010000: out_v[170] = 10'b0001010101;
    16'b0001000010010000: out_v[170] = 10'b0100010101;
    16'b0001000001111010: out_v[170] = 10'b0101010000;
    16'b0001000001010010: out_v[170] = 10'b1111001001;
    16'b0001000000110010: out_v[170] = 10'b1001011001;
    16'b0000000111010001: out_v[170] = 10'b1110110010;
    16'b0001000001110010: out_v[170] = 10'b1011010111;
    16'b0001000111010010: out_v[170] = 10'b0010101111;
    16'b0001000111110000: out_v[170] = 10'b0011011011;
    16'b0000000111010000: out_v[170] = 10'b1101100110;
    16'b0000000101010011: out_v[170] = 10'b1011010111;
    16'b0001000101111010: out_v[170] = 10'b0011001111;
    16'b0000000100110010: out_v[170] = 10'b1011001111;
    16'b0001000001101010: out_v[170] = 10'b1001110011;
    16'b0001000111000001: out_v[170] = 10'b0000111001;
    16'b0001000101010010: out_v[170] = 10'b0101110011;
    16'b0001000001010000: out_v[170] = 10'b0101001110;
    16'b0001000111000000: out_v[170] = 10'b0100010011;
    16'b0000000111110010: out_v[170] = 10'b0111011011;
    16'b0000000111010010: out_v[170] = 10'b1011011110;
    16'b0000000111010011: out_v[170] = 10'b1001111111;
    16'b0000000101010010: out_v[170] = 10'b0111010111;
    16'b0001000111010001: out_v[170] = 10'b0110111010;
    16'b0001000000101010: out_v[170] = 10'b1001011011;
    16'b0001000001100010: out_v[170] = 10'b1110010101;
    16'b0001000011110010: out_v[170] = 10'b0011001001;
    16'b0001000011010010: out_v[170] = 10'b0000001110;
    16'b0000000101110010: out_v[170] = 10'b0110001010;
    16'b0001000101010000: out_v[170] = 10'b0001001100;
    16'b0001000111110010: out_v[170] = 10'b0011110111;
    16'b0001000101010011: out_v[170] = 10'b0111011101;
    16'b0001000011111010: out_v[170] = 10'b1000101011;
    16'b0001000011000000: out_v[170] = 10'b0110001011;
    16'b0000000010000000: out_v[170] = 10'b1011100101;
    16'b0001000011110000: out_v[170] = 10'b0001011011;
    16'b0001000000111010: out_v[170] = 10'b0101101010;
    16'b0001000110000000: out_v[170] = 10'b0101010011;
    16'b0001000111110011: out_v[170] = 10'b1111110100;
    16'b0001000111010011: out_v[170] = 10'b1111101110;
    16'b0000000101110011: out_v[170] = 10'b0011010011;
    16'b0000000101111010: out_v[170] = 10'b0111011111;
    16'b0001000100000001: out_v[170] = 10'b0110000101;
    16'b0000000000000000: out_v[170] = 10'b1101010111;
    16'b0001000100000000: out_v[170] = 10'b0111100110;
    16'b0000000100000001: out_v[170] = 10'b1111000010;
    16'b0000000100000000: out_v[170] = 10'b0000111100;
    16'b0001000000000000: out_v[170] = 10'b1010101010;
    16'b0001000110000001: out_v[170] = 10'b1101011110;
    16'b0000000000000001: out_v[170] = 10'b1000110011;
    16'b0001000000000001: out_v[170] = 10'b0010111100;
    16'b0001000000010000: out_v[170] = 10'b0010111010;
    16'b0001000010000001: out_v[170] = 10'b1001011001;
    16'b0001000010010010: out_v[170] = 10'b1001100111;
    16'b0001000010000011: out_v[170] = 10'b0110101101;
    16'b0000000000010000: out_v[170] = 10'b0110100111;
    16'b0001000011000010: out_v[170] = 10'b0110000101;
    16'b0001000010000010: out_v[170] = 10'b0010101111;
    16'b0001000100010000: out_v[170] = 10'b1010101110;
    16'b0001000010010001: out_v[170] = 10'b0111010000;
    16'b0001000001000000: out_v[170] = 10'b1011011110;
    16'b0001000010110010: out_v[170] = 10'b1001001111;
    16'b0001000110010000: out_v[170] = 10'b1100110011;
    16'b0001000010010011: out_v[170] = 10'b1111011010;
    16'b0000000010010000: out_v[170] = 10'b0011111001;
    16'b0001000010110000: out_v[170] = 10'b0101010100;
    16'b0001000011000011: out_v[170] = 10'b1111001000;
    16'b0101000010110000: out_v[170] = 10'b1010111110;
    16'b0001000000110000: out_v[170] = 10'b1100101101;
    16'b0000000100010000: out_v[170] = 10'b1001000010;
    16'b0000000110000000: out_v[170] = 10'b1000101000;
    16'b0000000110010000: out_v[170] = 10'b0010010001;
    16'b0000000110000001: out_v[170] = 10'b1100111001;
    16'b0000000110010001: out_v[170] = 10'b0010111101;
    16'b0000000101010000: out_v[170] = 10'b1010001010;
    16'b0000000110010010: out_v[170] = 10'b0010111010;
    16'b0000000100010001: out_v[170] = 10'b0011001111;
    16'b0000000010000010: out_v[170] = 10'b0011110011;
    16'b0000000010000001: out_v[170] = 10'b0100110101;
    16'b0000000010010010: out_v[170] = 10'b1101111010;
    16'b0000000000000010: out_v[170] = 10'b0111101100;
    16'b0000000011000000: out_v[170] = 10'b0110110000;
    16'b0000000010100010: out_v[170] = 10'b0110111101;
    16'b0000000010001010: out_v[170] = 10'b1001110011;
    16'b0000000011100010: out_v[170] = 10'b0110110110;
    16'b0000000011011010: out_v[170] = 10'b1000010010;
    16'b0000000011000010: out_v[170] = 10'b0110010100;
    16'b0000000010000100: out_v[170] = 10'b1000011011;
    16'b0000000010000011: out_v[170] = 10'b1100100111;
    16'b0000000011010010: out_v[170] = 10'b1101011011;
    16'b0000000011011110: out_v[170] = 10'b1011101111;
    16'b0000000010010011: out_v[170] = 10'b1110000011;
    16'b0000000011001010: out_v[170] = 10'b1001010100;
    16'b0000000010011010: out_v[170] = 10'b0101100011;
    16'b0000000010110010: out_v[170] = 10'b1100011010;
    16'b0000000010011110: out_v[170] = 10'b1101110111;
    16'b0001000000000010: out_v[170] = 10'b1000100010;
    16'b0001000000010001: out_v[170] = 10'b1010110100;
    16'b0000000110000010: out_v[170] = 10'b1001001010;
    16'b0001000100010001: out_v[170] = 10'b1111000110;
    16'b0001000011010001: out_v[170] = 10'b0001101111;
    16'b0000000011010000: out_v[170] = 10'b1011001000;
    16'b0101000001110010: out_v[170] = 10'b1010010011;
    16'b0101000011110010: out_v[170] = 10'b1111100010;
    16'b0001000011100000: out_v[170] = 10'b1111001110;
    16'b0001000011110011: out_v[170] = 10'b1000011110;
    16'b0000000101000000: out_v[170] = 10'b1010011001;
    16'b1000000000000000: out_v[170] = 10'b0000011111;
    16'b1000000010000000: out_v[170] = 10'b1110001010;
    16'b0000000000001000: out_v[170] = 10'b0110101101;
    16'b1000000000000010: out_v[170] = 10'b0110001010;
    16'b0000000001000010: out_v[170] = 10'b0110110111;
    16'b1000000000001000: out_v[170] = 10'b0110110011;
    16'b0000000001000000: out_v[170] = 10'b0110111010;
    16'b0000000001010000: out_v[170] = 10'b1110100010;
    16'b1000000001000000: out_v[170] = 10'b1000111111;
    16'b1000000001010000: out_v[170] = 10'b0110110101;
    16'b0000000001011000: out_v[170] = 10'b0100011010;
    16'b0001000101000000: out_v[170] = 10'b1010010111;
    16'b0000000001001000: out_v[170] = 10'b0111101101;
    16'b1000000001001000: out_v[170] = 10'b0101110011;
    16'b0000000111000000: out_v[170] = 10'b1100000110;
    16'b0000000010010100: out_v[170] = 10'b1000101010;
    16'b0001000001000010: out_v[170] = 10'b1001001010;
    16'b1000000010000010: out_v[170] = 10'b1101100110;
    default: out_v[170] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001000000000000: out_v[171] = 10'b1001001010;
    16'b1000000100100000: out_v[171] = 10'b1000010011;
    16'b1001000100100101: out_v[171] = 10'b0011100001;
    16'b1001000100100001: out_v[171] = 10'b1011011111;
    16'b1000000000100000: out_v[171] = 10'b0110001000;
    16'b0000000000000000: out_v[171] = 10'b1100001011;
    16'b0001000000100001: out_v[171] = 10'b1000111110;
    16'b0000000000100101: out_v[171] = 10'b1100011011;
    16'b1000000100000101: out_v[171] = 10'b0011011111;
    16'b1000000000000101: out_v[171] = 10'b0010010011;
    16'b1001000100000101: out_v[171] = 10'b1100010011;
    16'b0000000100000000: out_v[171] = 10'b0000110001;
    16'b1000000000100001: out_v[171] = 10'b1010101111;
    16'b1000000100100101: out_v[171] = 10'b0111100000;
    16'b0000000100100000: out_v[171] = 10'b0101100011;
    16'b1000000100100001: out_v[171] = 10'b1110011001;
    16'b0001000100100001: out_v[171] = 10'b1100110100;
    16'b1000000000000000: out_v[171] = 10'b0000101010;
    16'b1001000000100001: out_v[171] = 10'b0110011100;
    16'b0001000000000001: out_v[171] = 10'b1000010011;
    16'b1000000100000100: out_v[171] = 10'b1111001000;
    16'b1000000100000000: out_v[171] = 10'b1100100011;
    16'b1000000100000001: out_v[171] = 10'b0100011110;
    16'b1000100100100000: out_v[171] = 10'b1101000000;
    16'b1001000000100101: out_v[171] = 10'b1001110111;
    16'b1000000000000100: out_v[171] = 10'b0000001011;
    16'b1000100100100001: out_v[171] = 10'b1010110101;
    16'b0001000000100101: out_v[171] = 10'b0010010111;
    16'b0001000100000000: out_v[171] = 10'b1111101111;
    16'b1100000100100000: out_v[171] = 10'b1011101011;
    16'b1000000000100101: out_v[171] = 10'b0110111110;
    16'b1001000000000101: out_v[171] = 10'b0010010001;
    16'b1001000100000001: out_v[171] = 10'b1101100001;
    16'b0001000100000001: out_v[171] = 10'b1101010110;
    16'b0000000000100000: out_v[171] = 10'b1100100000;
    16'b0000000100100001: out_v[171] = 10'b0111101100;
    16'b0100000100000000: out_v[171] = 10'b0101001000;
    16'b0100000000000000: out_v[171] = 10'b1101010010;
    16'b0101000000000000: out_v[171] = 10'b1101000110;
    16'b1100000100000000: out_v[171] = 10'b1101010000;
    16'b1100000000000000: out_v[171] = 10'b1110001010;
    16'b0101000010000000: out_v[171] = 10'b0001111010;
    16'b0000000100000001: out_v[171] = 10'b0111011111;
    16'b0101000110000000: out_v[171] = 10'b1010010011;
    16'b0101000100000001: out_v[171] = 10'b1100011010;
    16'b0100000100000001: out_v[171] = 10'b1000000111;
    16'b0101000000000001: out_v[171] = 10'b0001111101;
    16'b0100000000000001: out_v[171] = 10'b0100011110;
    16'b1100000000100000: out_v[171] = 10'b1101000001;
    16'b0100000010000001: out_v[171] = 10'b1100010011;
    16'b0101000100000000: out_v[171] = 10'b1001010111;
    16'b1101000100000000: out_v[171] = 10'b1011110101;
    16'b1100000100000001: out_v[171] = 10'b0011000100;
    16'b0100000010000000: out_v[171] = 10'b1011100001;
    16'b1101000000100000: out_v[171] = 10'b1110000110;
    16'b0101000110000001: out_v[171] = 10'b0010101111;
    16'b0000000000000001: out_v[171] = 10'b1110001110;
    16'b0100010010000001: out_v[171] = 10'b1111110111;
    16'b0101010010000001: out_v[171] = 10'b1010101110;
    16'b1101000100100000: out_v[171] = 10'b0110011110;
    16'b0100000110000001: out_v[171] = 10'b0011100111;
    16'b0100000000000100: out_v[171] = 10'b0110110101;
    16'b1101000110000000: out_v[171] = 10'b0101100110;
    16'b1101100000000000: out_v[171] = 10'b0111111001;
    16'b0101010010000000: out_v[171] = 10'b0010011111;
    16'b0101000010000001: out_v[171] = 10'b1011010010;
    16'b0100010110000001: out_v[171] = 10'b0011101011;
    16'b1100000000000001: out_v[171] = 10'b0000110110;
    16'b1101000000000000: out_v[171] = 10'b0010110101;
    16'b1100000000100001: out_v[171] = 10'b1110001110;
    16'b1100100100100000: out_v[171] = 10'b0011011001;
    16'b1100000100100001: out_v[171] = 10'b1010110110;
    16'b0001000010000001: out_v[171] = 10'b1000101001;
    16'b1010100100000000: out_v[171] = 10'b1100011100;
    16'b0000000010000000: out_v[171] = 10'b1100110010;
    16'b1000100100000000: out_v[171] = 10'b0101011010;
    16'b0001000110000001: out_v[171] = 10'b0111111000;
    16'b0000100100000000: out_v[171] = 10'b1011100101;
    16'b0001000010000000: out_v[171] = 10'b1001111100;
    16'b0001000110000000: out_v[171] = 10'b0101010110;
    16'b1010000100000000: out_v[171] = 10'b1111010111;
    16'b0000000110000000: out_v[171] = 10'b1111101110;
    16'b1001000110000001: out_v[171] = 10'b0100001000;
    16'b0001010010000001: out_v[171] = 10'b1000001011;
    16'b0001010110000001: out_v[171] = 10'b0011101101;
    16'b1100100100000000: out_v[171] = 10'b1011110101;
    16'b0100000000100000: out_v[171] = 10'b1101101010;
    16'b1100000000000100: out_v[171] = 10'b1010011110;
    16'b1001000000000001: out_v[171] = 10'b0001111011;
    16'b1001000100000000: out_v[171] = 10'b0011100110;
    16'b1001000000000000: out_v[171] = 10'b0001111000;
    16'b0100000000100101: out_v[171] = 10'b1011111011;
    16'b0100000000100001: out_v[171] = 10'b1100101110;
    16'b0100000000000101: out_v[171] = 10'b0111100110;
    16'b0100000000100100: out_v[171] = 10'b1101101010;
    16'b0101000000100001: out_v[171] = 10'b1011001011;
    16'b1100000000000010: out_v[171] = 10'b1101001001;
    16'b1100000100100010: out_v[171] = 10'b1001000011;
    16'b1100000100000010: out_v[171] = 10'b1111001001;
    16'b1100000000100010: out_v[171] = 10'b1001101111;
    16'b0100000100100000: out_v[171] = 10'b1110011000;
    default: out_v[171] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100000010010001: out_v[172] = 10'b1000001011;
    16'b0100000011010001: out_v[172] = 10'b1000110011;
    16'b0100100011010000: out_v[172] = 10'b1111011110;
    16'b0100100010010000: out_v[172] = 10'b1111001110;
    16'b0000000011010001: out_v[172] = 10'b1111110010;
    16'b0000000011010000: out_v[172] = 10'b0110111000;
    16'b0100000011110000: out_v[172] = 10'b0010001111;
    16'b0000000001010000: out_v[172] = 10'b0110110011;
    16'b0000000010000000: out_v[172] = 10'b1011001001;
    16'b0100100010000000: out_v[172] = 10'b1100100011;
    16'b0000000010000001: out_v[172] = 10'b0001110101;
    16'b0100000011000000: out_v[172] = 10'b1001101101;
    16'b0100000011010101: out_v[172] = 10'b0110001101;
    16'b0100100010010001: out_v[172] = 10'b1101011100;
    16'b0000000010010001: out_v[172] = 10'b1110001011;
    16'b0000100010010001: out_v[172] = 10'b1110110011;
    16'b0000000010010000: out_v[172] = 10'b0010010110;
    16'b0100000011010000: out_v[172] = 10'b1110000001;
    16'b0100000010010000: out_v[172] = 10'b1000000111;
    16'b0100100010110000: out_v[172] = 10'b0111101001;
    16'b0100000010000000: out_v[172] = 10'b1101001000;
    16'b0000000011000001: out_v[172] = 10'b1111001101;
    16'b0100100011010001: out_v[172] = 10'b0001010111;
    16'b0100000011000001: out_v[172] = 10'b1101100100;
    16'b0000100010000000: out_v[172] = 10'b0000000101;
    16'b0100100110010000: out_v[172] = 10'b1011001110;
    16'b0000100011010001: out_v[172] = 10'b0011110000;
    16'b0000100010010000: out_v[172] = 10'b1011000101;
    16'b0100000010110000: out_v[172] = 10'b1011101011;
    16'b0100000010000001: out_v[172] = 10'b1001001010;
    16'b0100000010010101: out_v[172] = 10'b0110010111;
    16'b0100000001010101: out_v[172] = 10'b1111000111;
    16'b0000100011010000: out_v[172] = 10'b0100110010;
    16'b0000000011000100: out_v[172] = 10'b1001010011;
    16'b0100000011000100: out_v[172] = 10'b1110100001;
    16'b0000000001000100: out_v[172] = 10'b0110000110;
    16'b0000000011000000: out_v[172] = 10'b1000011110;
    16'b0000000001000000: out_v[172] = 10'b0110001010;
    16'b0100000001000100: out_v[172] = 10'b1111101001;
    16'b0000100000000100: out_v[172] = 10'b1101001011;
    16'b0000000000000100: out_v[172] = 10'b0011011101;
    16'b0000000000000000: out_v[172] = 10'b0011010011;
    16'b0000100001000100: out_v[172] = 10'b1110000001;
    16'b0100000001000000: out_v[172] = 10'b0101111010;
    16'b0000000001000101: out_v[172] = 10'b0100010101;
    16'b0000000011000101: out_v[172] = 10'b1101010111;
    16'b0000100011000100: out_v[172] = 10'b1001111111;
    16'b0000100111000100: out_v[172] = 10'b0011010101;
    16'b0000100010010101: out_v[172] = 10'b0110000110;
    16'b0000100110000100: out_v[172] = 10'b1111011111;
    16'b0000000010000100: out_v[172] = 10'b0110100001;
    16'b0000100101000100: out_v[172] = 10'b0100011100;
    16'b0000100011000000: out_v[172] = 10'b0101010000;
    16'b0000100001000000: out_v[172] = 10'b1000011101;
    16'b0000100010000100: out_v[172] = 10'b0001100110;
    16'b0000000000000101: out_v[172] = 10'b1000000100;
    16'b0100000010010100: out_v[172] = 10'b0011111100;
    16'b0100100010010100: out_v[172] = 10'b0001001010;
    16'b0000100010000101: out_v[172] = 10'b0010110110;
    16'b0100100100010100: out_v[172] = 10'b1110001011;
    16'b0100000000010101: out_v[172] = 10'b1111000010;
    16'b0100000000010100: out_v[172] = 10'b1000110011;
    16'b0000000000010100: out_v[172] = 10'b1001000110;
    16'b0000100000000101: out_v[172] = 10'b1000001111;
    16'b0000100011000101: out_v[172] = 10'b1010001001;
    16'b0000100000010100: out_v[172] = 10'b0100001110;
    16'b0100100010010101: out_v[172] = 10'b1001001010;
    16'b0100100000010100: out_v[172] = 10'b0100111011;
    16'b0000100001000101: out_v[172] = 10'b1001011100;
    16'b0000100010010100: out_v[172] = 10'b0101011001;
    16'b0100000000000100: out_v[172] = 10'b1000010100;
    16'b0000100111000000: out_v[172] = 10'b1011110111;
    16'b0100100000010101: out_v[172] = 10'b0010011010;
    16'b0000000010000101: out_v[172] = 10'b1101100110;
    16'b0000100100000100: out_v[172] = 10'b0111000010;
    16'b0000100101000000: out_v[172] = 10'b0110011011;
    16'b0000000010010100: out_v[172] = 10'b1001011100;
    16'b0100100110010100: out_v[172] = 10'b1100111100;
    16'b0100000001010100: out_v[172] = 10'b0010001110;
    16'b0000000000010101: out_v[172] = 10'b1101000111;
    16'b0100000011010100: out_v[172] = 10'b1100010110;
    16'b0000100011000001: out_v[172] = 10'b0100001001;
    16'b0100100011000000: out_v[172] = 10'b0101101011;
    16'b0010100011000101: out_v[172] = 10'b0011001110;
    16'b0000100001000001: out_v[172] = 10'b1010000101;
    16'b0010100011000001: out_v[172] = 10'b1101100110;
    16'b0100100011000001: out_v[172] = 10'b0111001010;
    16'b0100100011010101: out_v[172] = 10'b0010110011;
    16'b0100100011010100: out_v[172] = 10'b0101100011;
    16'b0000100010000001: out_v[172] = 10'b0000110110;
    16'b0100100011000101: out_v[172] = 10'b1010100110;
    16'b0100000011000101: out_v[172] = 10'b1001110011;
    16'b0100100011000100: out_v[172] = 10'b1011000011;
    16'b0010100011000000: out_v[172] = 10'b1111111111;
    16'b0000000011010101: out_v[172] = 10'b0011110010;
    16'b0000100000000001: out_v[172] = 10'b0011010111;
    16'b0000000010010101: out_v[172] = 10'b1101000000;
    16'b0100000010000101: out_v[172] = 10'b0101011010;
    16'b0000000000000001: out_v[172] = 10'b0011100001;
    16'b0100000000000101: out_v[172] = 10'b0001110110;
    16'b0000100000010101: out_v[172] = 10'b1101001101;
    16'b0100100000010001: out_v[172] = 10'b1000011010;
    16'b0100000000010001: out_v[172] = 10'b0100011010;
    16'b0100000000110101: out_v[172] = 10'b0001110111;
    16'b0100000000110100: out_v[172] = 10'b1001110000;
    16'b0100100000000101: out_v[172] = 10'b1010100111;
    16'b0100100010000001: out_v[172] = 10'b1000110011;
    16'b0100100010000101: out_v[172] = 10'b1110110000;
    16'b0100000010000100: out_v[172] = 10'b0111011000;
    16'b0100000001000001: out_v[172] = 10'b0100100110;
    16'b0100000000000001: out_v[172] = 10'b0000111011;
    16'b0100000001000101: out_v[172] = 10'b1110100110;
    16'b0000000001010101: out_v[172] = 10'b1001100001;
    16'b0000100110000001: out_v[172] = 10'b0011110010;
    16'b0000000001000001: out_v[172] = 10'b1100000011;
    16'b0000100000010000: out_v[172] = 10'b1001011011;
    16'b0000000000010001: out_v[172] = 10'b1010111011;
    16'b0000100000010001: out_v[172] = 10'b0001011111;
    16'b0000100001010001: out_v[172] = 10'b0001001110;
    16'b0000000001010100: out_v[172] = 10'b1100101101;
    16'b0000000011010100: out_v[172] = 10'b1110101001;
    16'b0100000011110100: out_v[172] = 10'b0011101110;
    16'b0000100011010100: out_v[172] = 10'b0011111111;
    16'b0000000001110000: out_v[172] = 10'b0110111111;
    16'b0100000001010000: out_v[172] = 10'b0010001100;
    16'b0000000000010000: out_v[172] = 10'b1111101100;
    16'b0000000001010001: out_v[172] = 10'b1111100011;
    16'b0100000001110000: out_v[172] = 10'b0111001010;
    16'b0000100011010101: out_v[172] = 10'b0110100010;
    16'b0100100010000100: out_v[172] = 10'b1100110111;
    16'b0000100001010101: out_v[172] = 10'b0010110011;
    default: out_v[172] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000000100000: out_v[173] = 10'b1001001001;
    16'b0010000011110100: out_v[173] = 10'b0100011101;
    16'b0010100011010100: out_v[173] = 10'b1110011110;
    16'b0010100000000100: out_v[173] = 10'b0101010110;
    16'b1010100000000100: out_v[173] = 10'b0101101011;
    16'b0010000010000100: out_v[173] = 10'b1001001111;
    16'b0010100001000100: out_v[173] = 10'b1001000111;
    16'b0010100011000100: out_v[173] = 10'b1010000011;
    16'b1010100001000100: out_v[173] = 10'b1000010011;
    16'b0010000010100100: out_v[173] = 10'b1100010100;
    16'b0010000011000100: out_v[173] = 10'b0110011100;
    16'b1010000000100100: out_v[173] = 10'b0101010011;
    16'b0010000011100100: out_v[173] = 10'b0110100101;
    16'b0000000000110000: out_v[173] = 10'b1000101001;
    16'b0000000000000000: out_v[173] = 10'b1110001001;
    16'b1000000000110000: out_v[173] = 10'b0000101101;
    16'b0010000000100100: out_v[173] = 10'b0000010110;
    16'b0000000010100000: out_v[173] = 10'b0011111000;
    16'b0010000000010100: out_v[173] = 10'b1001010011;
    16'b0010100000010100: out_v[173] = 10'b1010011101;
    16'b0010100000100100: out_v[173] = 10'b0101110000;
    16'b0010000000000100: out_v[173] = 10'b1000101111;
    16'b0000100000000000: out_v[173] = 10'b0110101110;
    16'b1010000010100100: out_v[173] = 10'b0101000110;
    16'b0010100011110100: out_v[173] = 10'b1111011101;
    16'b1010000011100100: out_v[173] = 10'b1110010001;
    16'b0010000011010100: out_v[173] = 10'b0011101111;
    16'b0000100000100000: out_v[173] = 10'b0111010110;
    16'b0010100011100100: out_v[173] = 10'b1110110010;
    16'b1000000000100000: out_v[173] = 10'b0111010011;
    16'b1010100011000100: out_v[173] = 10'b0111011110;
    16'b1010000011000100: out_v[173] = 10'b1111100111;
    16'b0010000000110100: out_v[173] = 10'b0111110011;
    16'b0000000000010000: out_v[173] = 10'b0111100100;
    16'b0010000010110100: out_v[173] = 10'b0110110110;
    16'b1010100011010100: out_v[173] = 10'b0001110011;
    16'b1010100011100100: out_v[173] = 10'b1000110111;
    16'b0010000000100000: out_v[173] = 10'b0010010001;
    16'b1000000000000000: out_v[173] = 10'b1110001010;
    16'b1000000000010000: out_v[173] = 10'b1111011100;
    16'b1000000010000000: out_v[173] = 10'b0100110010;
    16'b1100000000000000: out_v[173] = 10'b0110001101;
    16'b0110000000100100: out_v[173] = 10'b0100011110;
    16'b0100000000000000: out_v[173] = 10'b1101001111;
    16'b0010000000000000: out_v[173] = 10'b0011001100;
    16'b0100000000100000: out_v[173] = 10'b0010100110;
    16'b1000000000000010: out_v[173] = 10'b0110010100;
    16'b1010100000100100: out_v[173] = 10'b1100001110;
    16'b1100000000100000: out_v[173] = 10'b1001001101;
    16'b0110000000000100: out_v[173] = 10'b1001110101;
    16'b0000000000000010: out_v[173] = 10'b1011001010;
    16'b1110000000100100: out_v[173] = 10'b1001010110;
    16'b1010000000000100: out_v[173] = 10'b1010111010;
    16'b1000100000000000: out_v[173] = 10'b1010101100;
    16'b1000100000100000: out_v[173] = 10'b0100011101;
    16'b0000000010000000: out_v[173] = 10'b1010000011;
    16'b1010000010000100: out_v[173] = 10'b1000101010;
    16'b1010000000010100: out_v[173] = 10'b0001111101;
    16'b1000000000010010: out_v[173] = 10'b0110011111;
    16'b1000000000110010: out_v[173] = 10'b1011111110;
    16'b1000100000000010: out_v[173] = 10'b0011111110;
    16'b1110000000000100: out_v[173] = 10'b1001101000;
    16'b1010000010010100: out_v[173] = 10'b1010111110;
    16'b1000000010010000: out_v[173] = 10'b1001110000;
    16'b0000000000010010: out_v[173] = 10'b1110000100;
    16'b1010000000000000: out_v[173] = 10'b1001011010;
    16'b0000000010010000: out_v[173] = 10'b0111100000;
    16'b0000000010110000: out_v[173] = 10'b0000111011;
    16'b0000000000100010: out_v[173] = 10'b1100011111;
    16'b1010000001000100: out_v[173] = 10'b1010110010;
    16'b1000000010110000: out_v[173] = 10'b0101000100;
    16'b0010000010010100: out_v[173] = 10'b1010100001;
    16'b1000000010100000: out_v[173] = 10'b0100100111;
    16'b0010000010000000: out_v[173] = 10'b1100000111;
    16'b0100100000100000: out_v[173] = 10'b0010110110;
    16'b0010100000100000: out_v[173] = 10'b1011111010;
    16'b1100100000100000: out_v[173] = 10'b0110101111;
    16'b1000000011010000: out_v[173] = 10'b0011001011;
    16'b0000000010010010: out_v[173] = 10'b0101111111;
    16'b1000000000100010: out_v[173] = 10'b1110010100;
    16'b0000000001000000: out_v[173] = 10'b0111010010;
    16'b1010000010110100: out_v[173] = 10'b0111110110;
    16'b0000000001010000: out_v[173] = 10'b0010110010;
    16'b0000000011010000: out_v[173] = 10'b1011001010;
    default: out_v[173] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000100000000110: out_v[174] = 10'b1101110111;
    16'b0100100001000100: out_v[174] = 10'b1101010111;
    16'b1000101001001101: out_v[174] = 10'b1011111011;
    16'b0000100000000100: out_v[174] = 10'b0000111000;
    16'b1000001000001001: out_v[174] = 10'b0000000001;
    16'b0000101001000100: out_v[174] = 10'b1111001101;
    16'b1000001000001000: out_v[174] = 10'b0100011011;
    16'b1000101001001000: out_v[174] = 10'b1110001101;
    16'b0000101001001100: out_v[174] = 10'b0100100111;
    16'b0000100001000100: out_v[174] = 10'b1001000101;
    16'b0000100001001100: out_v[174] = 10'b0011010101;
    16'b0000000000000100: out_v[174] = 10'b1001001001;
    16'b1000101001001100: out_v[174] = 10'b1010110111;
    16'b0000101000000100: out_v[174] = 10'b0000111011;
    16'b0100100000000100: out_v[174] = 10'b0000101001;
    16'b0000101000001101: out_v[174] = 10'b0010111100;
    16'b1000101000001000: out_v[174] = 10'b1111111001;
    16'b1000101001001001: out_v[174] = 10'b1000011001;
    16'b0000101000000101: out_v[174] = 10'b1000100011;
    16'b0000100000000000: out_v[174] = 10'b1010110101;
    16'b0000101001001101: out_v[174] = 10'b0000111011;
    16'b0100100001001100: out_v[174] = 10'b1011001000;
    16'b0100101001000100: out_v[174] = 10'b0001111001;
    16'b0000101000001001: out_v[174] = 10'b1101111110;
    16'b1000101000001001: out_v[174] = 10'b0001110011;
    16'b0100101001001100: out_v[174] = 10'b0110111000;
    16'b0000101001001000: out_v[174] = 10'b1111010111;
    16'b0000101000001100: out_v[174] = 10'b1111101010;
    16'b0100101000000100: out_v[174] = 10'b1010011010;
    16'b0000101000000111: out_v[174] = 10'b0011011111;
    16'b0000100000001100: out_v[174] = 10'b1110111011;
    16'b0000101000001000: out_v[174] = 10'b1011110011;
    16'b0000000000000000: out_v[174] = 10'b0011110000;
    16'b0000101001001001: out_v[174] = 10'b1010011111;
    16'b0000100000000010: out_v[174] = 10'b0001011100;
    16'b0000101000000000: out_v[174] = 10'b0001001110;
    16'b0000110000000000: out_v[174] = 10'b1110000010;
    16'b0000010000000010: out_v[174] = 10'b0101101011;
    16'b0000010000000000: out_v[174] = 10'b1100000011;
    16'b0100110000000000: out_v[174] = 10'b0100001001;
    16'b0000110000000010: out_v[174] = 10'b1111010010;
    16'b0100010000000000: out_v[174] = 10'b1000100011;
    16'b0000110000000100: out_v[174] = 10'b1111001010;
    16'b0000000000000001: out_v[174] = 10'b0100010111;
    16'b0000010000000100: out_v[174] = 10'b0011011001;
    16'b0000010000000001: out_v[174] = 10'b0000010101;
    16'b0000111000000100: out_v[174] = 10'b0010101110;
    16'b0000100000000101: out_v[174] = 10'b1011110010;
    16'b0100110000000100: out_v[174] = 10'b1101010000;
    16'b0100100000000000: out_v[174] = 10'b0010100101;
    16'b0000110000000001: out_v[174] = 10'b1011001110;
    16'b0000111000000000: out_v[174] = 10'b1100000110;
    16'b0000010000000101: out_v[174] = 10'b0001101010;
    16'b0000100000000001: out_v[174] = 10'b0101010011;
    16'b0000000000000101: out_v[174] = 10'b1110100100;
    16'b0000110000000101: out_v[174] = 10'b0110001011;
    16'b0100110000000001: out_v[174] = 10'b1001101110;
    16'b1000010000000100: out_v[174] = 10'b0100110101;
    16'b1000000000000100: out_v[174] = 10'b0100011110;
    16'b1000010000000101: out_v[174] = 10'b0110100101;
    16'b0100010000000100: out_v[174] = 10'b0010010011;
    16'b0000010000000110: out_v[174] = 10'b1010010111;
    16'b0000110000000110: out_v[174] = 10'b1110100100;
    16'b0100110000000111: out_v[174] = 10'b0011111111;
    16'b0000010000010111: out_v[174] = 10'b0000001111;
    16'b0000110000000111: out_v[174] = 10'b0101111011;
    16'b0000000000000110: out_v[174] = 10'b0011111111;
    16'b0100110000000110: out_v[174] = 10'b1010011101;
    16'b0000010000000111: out_v[174] = 10'b1001011000;
    16'b0100110000000101: out_v[174] = 10'b0100011001;
    16'b0000011001000000: out_v[174] = 10'b1000100100;
    16'b0000010001000000: out_v[174] = 10'b1100000000;
    16'b0000011001000100: out_v[174] = 10'b0000101101;
    16'b0000111000000001: out_v[174] = 10'b1110100010;
    16'b0000011000000000: out_v[174] = 10'b1001011011;
    16'b0000011000000100: out_v[174] = 10'b0110011111;
    16'b0000011000000101: out_v[174] = 10'b1101001001;
    16'b0000111000000101: out_v[174] = 10'b0100110000;
    16'b0000001000000101: out_v[174] = 10'b1110000011;
    16'b0000001000000000: out_v[174] = 10'b1111001000;
    16'b0000110000010010: out_v[174] = 10'b1011100111;
    16'b0000001001000100: out_v[174] = 10'b0111010010;
    16'b0000001001000101: out_v[174] = 10'b0110010000;
    16'b0000001000000100: out_v[174] = 10'b1101000110;
    16'b0000111000000110: out_v[174] = 10'b0011111000;
    16'b0000000001000100: out_v[174] = 10'b1000110110;
    16'b0000010000010010: out_v[174] = 10'b1000010110;
    16'b0000010001000100: out_v[174] = 10'b0001111010;
    16'b0000100000000111: out_v[174] = 10'b1001100101;
    16'b0000000001000000: out_v[174] = 10'b1000110110;
    16'b0000110001000000: out_v[174] = 10'b1110001000;
    16'b0000111000000111: out_v[174] = 10'b1111110111;
    16'b0000000010000000: out_v[174] = 10'b1010000111;
    16'b0000010010000100: out_v[174] = 10'b1011001101;
    16'b0000010000001100: out_v[174] = 10'b0000110110;
    16'b1000011000001001: out_v[174] = 10'b0011001010;
    16'b0000000010000100: out_v[174] = 10'b1101100110;
    16'b0000010010000000: out_v[174] = 10'b1000101101;
    16'b0000000001000101: out_v[174] = 10'b0011110011;
    16'b0000000000010111: out_v[174] = 10'b0111001010;
    16'b0000000000010011: out_v[174] = 10'b1100011010;
    16'b0000000000010101: out_v[174] = 10'b1111000111;
    16'b0000000000010010: out_v[174] = 10'b0111001111;
    16'b0010001000000101: out_v[174] = 10'b0111000111;
    16'b0000010000010011: out_v[174] = 10'b1011111111;
    16'b0000001001000000: out_v[174] = 10'b1100001101;
    16'b0000001000010111: out_v[174] = 10'b0101111101;
    16'b0000000000000010: out_v[174] = 10'b0100001101;
    16'b0000000000000011: out_v[174] = 10'b1001001101;
    16'b0000000000000111: out_v[174] = 10'b1100011111;
    16'b0010000000000101: out_v[174] = 10'b1111100110;
    16'b0000000000010001: out_v[174] = 10'b1101111010;
    16'b0000001000010110: out_v[174] = 10'b0110111111;
    16'b0000000001000001: out_v[174] = 10'b0011010011;
    16'b0000000000010000: out_v[174] = 10'b0111101111;
    16'b0000000000010110: out_v[174] = 10'b0111000110;
    16'b0100110001000000: out_v[174] = 10'b0010001010;
    16'b0000110000000011: out_v[174] = 10'b0100100100;
    16'b0000110000010011: out_v[174] = 10'b0101010101;
    16'b0000110001000011: out_v[174] = 10'b1011110111;
    16'b0000110001000010: out_v[174] = 10'b1011111010;
    16'b0000100000010010: out_v[174] = 10'b0110110000;
    16'b0000010000010000: out_v[174] = 10'b0110101001;
    16'b0000011000010110: out_v[174] = 10'b1101101011;
    16'b0000011000000001: out_v[174] = 10'b0001110011;
    16'b0000010000010110: out_v[174] = 10'b0000001111;
    16'b0010011000000101: out_v[174] = 10'b1000111001;
    16'b0000110000010110: out_v[174] = 10'b1101000110;
    16'b0000011000010010: out_v[174] = 10'b1111100101;
    default: out_v[174] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0110000011011000: out_v[175] = 10'b0011100100;
    16'b1000010001011000: out_v[175] = 10'b0111110001;
    16'b1010010011011000: out_v[175] = 10'b0011100110;
    16'b0010010011011000: out_v[175] = 10'b1011000101;
    16'b0000010001011000: out_v[175] = 10'b1011011011;
    16'b0010000001011000: out_v[175] = 10'b1100010111;
    16'b0010010001011000: out_v[175] = 10'b1111100011;
    16'b1010000000001000: out_v[175] = 10'b0000100111;
    16'b0111010011010000: out_v[175] = 10'b1110001011;
    16'b1010010001011000: out_v[175] = 10'b1010101011;
    16'b0000000001011000: out_v[175] = 10'b1011110001;
    16'b0010000011011000: out_v[175] = 10'b1111110110;
    16'b0111000011010000: out_v[175] = 10'b0010110000;
    16'b0110000011010000: out_v[175] = 10'b1011100011;
    16'b0011010011011000: out_v[175] = 10'b0111110111;
    16'b0110010011011000: out_v[175] = 10'b0010111001;
    16'b0011010001011000: out_v[175] = 10'b0000111011;
    16'b0010000000001000: out_v[175] = 10'b0001101011;
    16'b1000000001011000: out_v[175] = 10'b0011101101;
    16'b0011000011011000: out_v[175] = 10'b1010110001;
    16'b1000010000011000: out_v[175] = 10'b0011110101;
    16'b0110000010010000: out_v[175] = 10'b0101110000;
    16'b1010000001011000: out_v[175] = 10'b1010001010;
    16'b0010010010010000: out_v[175] = 10'b1010111111;
    16'b0111000011011000: out_v[175] = 10'b0011111101;
    16'b1000010000000000: out_v[175] = 10'b0100110011;
    16'b1010010000001000: out_v[175] = 10'b0011011111;
    16'b0010010000001000: out_v[175] = 10'b0010011001;
    16'b1000010000001000: out_v[175] = 10'b0111100110;
    16'b0110010011010000: out_v[175] = 10'b1011010101;
    16'b0110010010010000: out_v[175] = 10'b0111000010;
    16'b1110010011011000: out_v[175] = 10'b1100110001;
    16'b1000000000001000: out_v[175] = 10'b1000000100;
    16'b1010000011011000: out_v[175] = 10'b1110001010;
    16'b0111010011011000: out_v[175] = 10'b0011110011;
    16'b0011000001011000: out_v[175] = 10'b1001100100;
    16'b0010000010010000: out_v[175] = 10'b1100000010;
    16'b0010000011010000: out_v[175] = 10'b0001011011;
    16'b0111000010010000: out_v[175] = 10'b0111100011;
    16'b0010010011010000: out_v[175] = 10'b1110101011;
    16'b0000010000000000: out_v[175] = 10'b1011011010;
    16'b0000000000000000: out_v[175] = 10'b0010010111;
    16'b1000000000010000: out_v[175] = 10'b1011001010;
    16'b1000000001010000: out_v[175] = 10'b0010100110;
    16'b1000000000000000: out_v[175] = 10'b1011001001;
    16'b1001000011011000: out_v[175] = 10'b1100101011;
    16'b1001000001010000: out_v[175] = 10'b0011110011;
    16'b1000000011010000: out_v[175] = 10'b1011101011;
    16'b1000000011011000: out_v[175] = 10'b0011010011;
    16'b1001000011010000: out_v[175] = 10'b0111011000;
    16'b0000000000010000: out_v[175] = 10'b1111010001;
    16'b1001000001011000: out_v[175] = 10'b1100011010;
    16'b1001000000010000: out_v[175] = 10'b0011011111;
    16'b0001000001011000: out_v[175] = 10'b1011010100;
    16'b0101000011010000: out_v[175] = 10'b1010110111;
    16'b0101000011011000: out_v[175] = 10'b0110001001;
    16'b0001000000000000: out_v[175] = 10'b1010110101;
    16'b0000010000001000: out_v[175] = 10'b1010011110;
    16'b0100000011010000: out_v[175] = 10'b1000110101;
    16'b0001000000001000: out_v[175] = 10'b1001100000;
    16'b0001010000000000: out_v[175] = 10'b1011111111;
    16'b0010000000000000: out_v[175] = 10'b1001010110;
    16'b0101010011011000: out_v[175] = 10'b0010111010;
    16'b0001000000011000: out_v[175] = 10'b0011100111;
    16'b0100010010001000: out_v[175] = 10'b0001110111;
    16'b0001000000010000: out_v[175] = 10'b1001011110;
    16'b0001010000001000: out_v[175] = 10'b1000000111;
    16'b1001000000001000: out_v[175] = 10'b0100001110;
    16'b0001000011011000: out_v[175] = 10'b0010101111;
    16'b0000000000001000: out_v[175] = 10'b0011000100;
    16'b0001000100001000: out_v[175] = 10'b0111100110;
    16'b0001000001001000: out_v[175] = 10'b1001100110;
    16'b0011000000001000: out_v[175] = 10'b1111100010;
    16'b0001010001011000: out_v[175] = 10'b1001111110;
    16'b1010000000000000: out_v[175] = 10'b1010000101;
    16'b0001000011010000: out_v[175] = 10'b1010110100;
    16'b0100010011010000: out_v[175] = 10'b0000110101;
    16'b0010010000000000: out_v[175] = 10'b1000110010;
    16'b0101010011010000: out_v[175] = 10'b1111101011;
    16'b0000000010011000: out_v[175] = 10'b0000100101;
    16'b0100000010011000: out_v[175] = 10'b1100101001;
    16'b1100000011011000: out_v[175] = 10'b0000001010;
    16'b0100000010010000: out_v[175] = 10'b0101101101;
    16'b0100010010010000: out_v[175] = 10'b1100100101;
    16'b1000000010011000: out_v[175] = 10'b0101001100;
    16'b1100000011010000: out_v[175] = 10'b1011001010;
    16'b1100000010000000: out_v[175] = 10'b1010001010;
    16'b0100000010010010: out_v[175] = 10'b1000110100;
    16'b0100000010000000: out_v[175] = 10'b0001001111;
    16'b0000010011011000: out_v[175] = 10'b0000110101;
    16'b0000000010010000: out_v[175] = 10'b1111000101;
    16'b0000010000010000: out_v[175] = 10'b1100001111;
    16'b0000010000011000: out_v[175] = 10'b0100110110;
    16'b0100000011011000: out_v[175] = 10'b1011110011;
    16'b0001010011011000: out_v[175] = 10'b0000111011;
    16'b1100000010010000: out_v[175] = 10'b1111011100;
    16'b1100000010011000: out_v[175] = 10'b0101011001;
    16'b1101000010010000: out_v[175] = 10'b1111001111;
    16'b0101000010010000: out_v[175] = 10'b1000110111;
    16'b1101000011011000: out_v[175] = 10'b1110111010;
    16'b1000010011011000: out_v[175] = 10'b1010101000;
    16'b0000000011011000: out_v[175] = 10'b1000100100;
    16'b1001010001011000: out_v[175] = 10'b0110011010;
    16'b1101000011010000: out_v[175] = 10'b1100011100;
    16'b0000010001010000: out_v[175] = 10'b0101001100;
    16'b0000000001010000: out_v[175] = 10'b1100111000;
    16'b1110000011011000: out_v[175] = 10'b0010101111;
    16'b0110000010001000: out_v[175] = 10'b0010100000;
    16'b0110000010001010: out_v[175] = 10'b0001010110;
    16'b0010010000010000: out_v[175] = 10'b1100110000;
    16'b0010000000010000: out_v[175] = 10'b1001110000;
    16'b0010000001010000: out_v[175] = 10'b0100101100;
    16'b0000000010001000: out_v[175] = 10'b1100010111;
    16'b0010010001010000: out_v[175] = 10'b1100000000;
    16'b0010000010001000: out_v[175] = 10'b1101011010;
    16'b0010000011001000: out_v[175] = 10'b1101111111;
    16'b0010000000000010: out_v[175] = 10'b1110100001;
    16'b0010010010001000: out_v[175] = 10'b0101110110;
    16'b0110010010001010: out_v[175] = 10'b1001011011;
    16'b0110000000001010: out_v[175] = 10'b0010011111;
    16'b0110010010001000: out_v[175] = 10'b1111100010;
    16'b0010010011001000: out_v[175] = 10'b0111111111;
    16'b0100000010001000: out_v[175] = 10'b0011111010;
    16'b0000000000000010: out_v[175] = 10'b0100111010;
    16'b0000100000100100: out_v[175] = 10'b0100101111;
    16'b1000100000100100: out_v[175] = 10'b1111011110;
    16'b0110010010000000: out_v[175] = 10'b1101100011;
    16'b1000010000010000: out_v[175] = 10'b1111110001;
    16'b1000000000100000: out_v[175] = 10'b0100010101;
    16'b1000100000000100: out_v[175] = 10'b1001101000;
    16'b0110010010010010: out_v[175] = 10'b1000110111;
    16'b0110010010011000: out_v[175] = 10'b1011001011;
    16'b0010010010011000: out_v[175] = 10'b0101001010;
    16'b1000010001010000: out_v[175] = 10'b0101110100;
    16'b0000000001001000: out_v[175] = 10'b1101001111;
    16'b0011000001001000: out_v[175] = 10'b1101101001;
    16'b1000000000011000: out_v[175] = 10'b0101110110;
    16'b1000000001001000: out_v[175] = 10'b0111100010;
    16'b0010000001001000: out_v[175] = 10'b0100110011;
    16'b0000000000011000: out_v[175] = 10'b1111001000;
    16'b0000000011010000: out_v[175] = 10'b0101011100;
    16'b0000000001000000: out_v[175] = 10'b1101011000;
    16'b0011000001000000: out_v[175] = 10'b1111011110;
    16'b1010000000010000: out_v[175] = 10'b1010101011;
    16'b1110000010001000: out_v[175] = 10'b1001000101;
    16'b1010000001010000: out_v[175] = 10'b1011010011;
    16'b1010000010001000: out_v[175] = 10'b0111000011;
    16'b1010010000000000: out_v[175] = 10'b0011110110;
    16'b0110000010011000: out_v[175] = 10'b0011001101;
    16'b0010000010011000: out_v[175] = 10'b0001111010;
    16'b0000010010011000: out_v[175] = 10'b1001011100;
    16'b1010000000000010: out_v[175] = 10'b1111100010;
    default: out_v[175] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010100000000000: out_v[176] = 10'b0010110100;
    16'b0010100000100000: out_v[176] = 10'b0110010001;
    16'b0010100000100001: out_v[176] = 10'b1100010000;
    16'b0010000000100001: out_v[176] = 10'b0101001101;
    16'b0000100000100000: out_v[176] = 10'b0001101000;
    16'b0000100000100001: out_v[176] = 10'b0010011110;
    16'b0000000000100000: out_v[176] = 10'b0001001111;
    16'b0010001000100001: out_v[176] = 10'b1110000111;
    16'b0010000000100000: out_v[176] = 10'b0001001111;
    16'b0010101000100001: out_v[176] = 10'b1101000111;
    16'b0000101000100001: out_v[176] = 10'b1010110110;
    16'b0000000000100001: out_v[176] = 10'b1001011100;
    16'b0010000000000001: out_v[176] = 10'b0000001111;
    16'b0000001000100001: out_v[176] = 10'b1010111000;
    16'b0010000000000000: out_v[176] = 10'b0001011010;
    16'b0000001000000001: out_v[176] = 10'b1101100011;
    16'b0010100000000001: out_v[176] = 10'b0011011000;
    16'b0010101000000001: out_v[176] = 10'b1000100010;
    16'b0000100000000000: out_v[176] = 10'b0001110001;
    16'b0010001000000001: out_v[176] = 10'b1000111101;
    16'b0000000000000000: out_v[176] = 10'b0011000110;
    16'b0000000000000001: out_v[176] = 10'b1101000001;
    16'b0010101000100000: out_v[176] = 10'b0011001101;
    16'b0000001000000000: out_v[176] = 10'b0100110100;
    16'b0000011000100000: out_v[176] = 10'b1101011011;
    16'b0000010000100000: out_v[176] = 10'b1000100101;
    16'b0010001000000000: out_v[176] = 10'b0100001010;
    16'b0000001000100000: out_v[176] = 10'b0111010110;
    16'b0000000001100000: out_v[176] = 10'b1110000101;
    16'b0010001000100000: out_v[176] = 10'b1111011101;
    16'b0000010000100001: out_v[176] = 10'b1000111010;
    16'b0000011000000000: out_v[176] = 10'b0101110001;
    16'b0000000001100001: out_v[176] = 10'b0001011010;
    16'b0010011000000001: out_v[176] = 10'b1000111011;
    16'b0000011000100001: out_v[176] = 10'b0011100111;
    16'b0000100000000001: out_v[176] = 10'b1011000100;
    16'b0000101000100000: out_v[176] = 10'b0011011001;
    16'b0000011000000001: out_v[176] = 10'b0001010101;
    16'b0010011000100001: out_v[176] = 10'b1010110101;
    16'b0010101000000000: out_v[176] = 10'b1011001111;
    16'b0010000000000011: out_v[176] = 10'b1101011111;
    16'b0000101000000001: out_v[176] = 10'b0110000011;
    16'b0000000000000011: out_v[176] = 10'b1101011011;
    16'b0000101000000000: out_v[176] = 10'b0011011011;
    16'b0010100000000010: out_v[176] = 10'b0110110100;
    16'b0010100000000011: out_v[176] = 10'b0010001011;
    16'b0000100000001001: out_v[176] = 10'b0110111010;
    16'b0000000000000101: out_v[176] = 10'b0001100101;
    16'b0000100000001000: out_v[176] = 10'b0110000001;
    16'b0000100000000101: out_v[176] = 10'b0010000001;
    16'b0000000000001001: out_v[176] = 10'b1001010101;
    16'b0010000000000010: out_v[176] = 10'b1011000100;
    16'b0010100000001001: out_v[176] = 10'b1101011111;
    16'b0010100000001011: out_v[176] = 10'b0111010011;
    16'b0000100000000100: out_v[176] = 10'b1110000110;
    16'b0000100000000010: out_v[176] = 10'b1101101010;
    16'b0000000000001000: out_v[176] = 10'b1101110011;
    16'b0000000000000100: out_v[176] = 10'b1101001111;
    default: out_v[176] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1000101110001010: out_v[177] = 10'b0010001101;
    16'b1000101110001000: out_v[177] = 10'b1100001011;
    16'b0000001100001010: out_v[177] = 10'b1001011100;
    16'b0010101100001010: out_v[177] = 10'b0111111110;
    16'b1000100110011000: out_v[177] = 10'b0010110011;
    16'b0000101000000010: out_v[177] = 10'b1000010111;
    16'b1010101000000010: out_v[177] = 10'b0100010111;
    16'b1000101110011010: out_v[177] = 10'b0101001011;
    16'b0000101110000000: out_v[177] = 10'b1111010111;
    16'b0000101100000000: out_v[177] = 10'b0100011001;
    16'b1000101110000010: out_v[177] = 10'b1111000111;
    16'b0000101100000010: out_v[177] = 10'b0110010011;
    16'b1000001110001010: out_v[177] = 10'b1000011001;
    16'b1010001110001010: out_v[177] = 10'b0010110111;
    16'b0000100110000000: out_v[177] = 10'b1111010011;
    16'b0000001100000010: out_v[177] = 10'b1000100100;
    16'b1010101110001010: out_v[177] = 10'b1111110011;
    16'b1010101100001010: out_v[177] = 10'b1011111101;
    16'b0000101100001010: out_v[177] = 10'b0110110001;
    16'b0010101110001010: out_v[177] = 10'b1011011011;
    16'b0010101000000010: out_v[177] = 10'b1111110100;
    16'b0001100110011000: out_v[177] = 10'b0101110110;
    16'b1010101010001010: out_v[177] = 10'b1110110010;
    16'b1000101010001010: out_v[177] = 10'b0110011010;
    16'b0000101110001010: out_v[177] = 10'b0101001001;
    16'b1000101100001010: out_v[177] = 10'b1001010111;
    16'b1010101000001010: out_v[177] = 10'b1011101111;
    16'b1000101110000000: out_v[177] = 10'b1011000011;
    16'b0000101110000010: out_v[177] = 10'b1011100110;
    16'b1000001100001010: out_v[177] = 10'b0000011111;
    16'b1001100110011000: out_v[177] = 10'b1001000111;
    16'b1000101110011000: out_v[177] = 10'b1100010011;
    16'b0000101010001010: out_v[177] = 10'b1000000011;
    16'b1000101000001010: out_v[177] = 10'b0001110110;
    16'b0010101100000010: out_v[177] = 10'b1110111110;
    16'b0000101110001000: out_v[177] = 10'b0010101111;
    16'b0000001110001010: out_v[177] = 10'b1001011010;
    16'b0010101000001010: out_v[177] = 10'b0000111011;
    16'b1010001010001010: out_v[177] = 10'b0110010001;
    16'b0000101000001010: out_v[177] = 10'b1110110010;
    16'b1000101100000010: out_v[177] = 10'b1010011111;
    16'b1000101000000010: out_v[177] = 10'b1100011111;
    16'b0010101010001010: out_v[177] = 10'b0110001011;
    16'b0000100100000010: out_v[177] = 10'b1110111011;
    16'b0001100110010000: out_v[177] = 10'b0101100101;
    16'b1001101110011010: out_v[177] = 10'b1010001110;
    16'b0001100000001000: out_v[177] = 10'b0101100111;
    16'b0001000100000000: out_v[177] = 10'b1101100110;
    16'b0000000100000000: out_v[177] = 10'b1001101011;
    16'b0011000100000000: out_v[177] = 10'b1111001110;
    16'b0001001100000000: out_v[177] = 10'b0001101011;
    16'b0000100000000000: out_v[177] = 10'b1101100001;
    16'b0010000100000000: out_v[177] = 10'b1110100101;
    16'b0011001100000000: out_v[177] = 10'b1010000011;
    16'b0000000000000000: out_v[177] = 10'b0000101111;
    16'b1000000000001000: out_v[177] = 10'b1000100011;
    16'b0000100100000000: out_v[177] = 10'b1110000111;
    16'b0001100100000000: out_v[177] = 10'b0000101111;
    16'b0001001000000000: out_v[177] = 10'b1011011101;
    16'b0001100000000000: out_v[177] = 10'b1001110001;
    16'b0011100100000000: out_v[177] = 10'b1010110011;
    16'b1000100000000000: out_v[177] = 10'b1110110011;
    16'b0000000000001000: out_v[177] = 10'b1011111100;
    16'b0001000000000000: out_v[177] = 10'b1110110001;
    16'b1000000000000000: out_v[177] = 10'b1101101001;
    16'b0010101000000000: out_v[177] = 10'b0110011101;
    16'b1011100000000000: out_v[177] = 10'b1110111111;
    16'b1010101000000000: out_v[177] = 10'b0010000100;
    16'b1011100010011000: out_v[177] = 10'b0010100010;
    16'b1011100000011000: out_v[177] = 10'b1011101011;
    16'b0011100010011000: out_v[177] = 10'b1001010111;
    16'b1011101010011010: out_v[177] = 10'b0010111111;
    16'b1011100010010000: out_v[177] = 10'b1110110110;
    16'b1001100010011000: out_v[177] = 10'b0101010110;
    16'b0011101010011000: out_v[177] = 10'b1000111010;
    16'b0011100010010000: out_v[177] = 10'b0110011111;
    16'b1011101000000000: out_v[177] = 10'b1110111011;
    16'b1011100010011010: out_v[177] = 10'b1111000011;
    16'b0011101000000000: out_v[177] = 10'b1011000110;
    16'b0010101000001000: out_v[177] = 10'b1001011100;
    16'b1011101010011000: out_v[177] = 10'b0011001011;
    16'b0011101000001000: out_v[177] = 10'b0100111000;
    16'b1011101000001000: out_v[177] = 10'b1111111011;
    16'b0001100010011000: out_v[177] = 10'b1111001101;
    16'b1001101110011000: out_v[177] = 10'b0010110011;
    16'b1010101000001000: out_v[177] = 10'b1011110111;
    16'b1001100110011010: out_v[177] = 10'b1001100110;
    16'b0000101010000010: out_v[177] = 10'b0110100001;
    16'b0000101000010000: out_v[177] = 10'b1110100111;
    16'b0010101010001000: out_v[177] = 10'b0000011011;
    16'b0000001000010000: out_v[177] = 10'b0011111011;
    16'b0000001110000000: out_v[177] = 10'b1100001011;
    16'b0000101010010000: out_v[177] = 10'b1010011111;
    16'b0000001010000000: out_v[177] = 10'b0111001111;
    16'b0010101000011000: out_v[177] = 10'b1011111011;
    16'b0001001100010000: out_v[177] = 10'b0111011110;
    16'b0000001100010010: out_v[177] = 10'b1110100011;
    16'b0000001111100000: out_v[177] = 10'b0110001011;
    16'b0010101010000000: out_v[177] = 10'b0001011100;
    16'b0000101010000000: out_v[177] = 10'b0011101010;
    16'b0000101010011000: out_v[177] = 10'b1111110100;
    16'b0000101010001000: out_v[177] = 10'b0101011011;
    16'b0010101010011000: out_v[177] = 10'b0000001111;
    16'b0000001100010000: out_v[177] = 10'b0001101000;
    16'b0010101000010000: out_v[177] = 10'b0001111011;
    16'b0010001110000000: out_v[177] = 10'b0000011111;
    16'b0000001110010000: out_v[177] = 10'b1110100101;
    16'b0000101000011000: out_v[177] = 10'b1111011111;
    16'b0000101110011010: out_v[177] = 10'b1000001011;
    16'b0000001111000000: out_v[177] = 10'b1100010011;
    16'b0000101000010010: out_v[177] = 10'b1010101011;
    16'b0000001110000010: out_v[177] = 10'b0000111010;
    16'b0010001000010000: out_v[177] = 10'b0111111001;
    16'b0010101110000000: out_v[177] = 10'b1111010110;
    16'b0010101010010000: out_v[177] = 10'b0111100110;
    16'b0010001010000000: out_v[177] = 10'b1001111101;
    16'b0000001110010010: out_v[177] = 10'b1101101111;
    16'b0001101010011010: out_v[177] = 10'b0101111110;
    16'b0001000010001000: out_v[177] = 10'b1111010100;
    16'b0001100000010000: out_v[177] = 10'b0010011111;
    16'b0001000000010010: out_v[177] = 10'b0100010111;
    16'b0001000000011010: out_v[177] = 10'b0010111011;
    16'b0001000010000010: out_v[177] = 10'b0111110011;
    16'b0001000010011010: out_v[177] = 10'b1000000111;
    16'b0001000010010010: out_v[177] = 10'b1001011100;
    16'b0001001010011000: out_v[177] = 10'b1101000111;
    16'b0001000010001010: out_v[177] = 10'b0010010111;
    16'b0001001010011010: out_v[177] = 10'b0011111111;
    16'b0001000000000010: out_v[177] = 10'b1001110001;
    16'b0001000000010000: out_v[177] = 10'b0111110001;
    16'b0001000000001010: out_v[177] = 10'b0010110111;
    16'b0001101000010010: out_v[177] = 10'b0101110011;
    16'b0001000000011000: out_v[177] = 10'b0101011010;
    16'b0001000110011010: out_v[177] = 10'b1001010011;
    16'b0001000010011000: out_v[177] = 10'b1111010011;
    16'b0000001010010010: out_v[177] = 10'b0101011010;
    16'b0000001010011010: out_v[177] = 10'b1011000100;
    16'b0001000110001000: out_v[177] = 10'b0011110110;
    16'b1001000010011010: out_v[177] = 10'b0110110011;
    16'b0001000100001000: out_v[177] = 10'b1001000000;
    16'b0001101000010000: out_v[177] = 10'b1111010011;
    16'b0000001010011000: out_v[177] = 10'b1011100001;
    16'b0000001000010010: out_v[177] = 10'b1101010011;
    16'b0001101010010000: out_v[177] = 10'b0101000110;
    16'b0001000000001000: out_v[177] = 10'b1011100010;
    16'b1001001010011010: out_v[177] = 10'b0001111010;
    16'b0001101010010010: out_v[177] = 10'b1111011111;
    16'b0001001000010010: out_v[177] = 10'b0000110011;
    16'b0001001010010010: out_v[177] = 10'b0100011010;
    16'b0001000110011000: out_v[177] = 10'b0011011010;
    16'b0000000010001000: out_v[177] = 10'b1010010001;
    16'b0001000010010000: out_v[177] = 10'b1011001111;
    16'b0001000010000000: out_v[177] = 10'b0101010011;
    16'b0001000110010000: out_v[177] = 10'b0100011000;
    16'b0001100010010010: out_v[177] = 10'b1101011010;
    16'b0001000100011000: out_v[177] = 10'b1001111011;
    16'b0001001000011010: out_v[177] = 10'b1110001111;
    16'b0001001000010000: out_v[177] = 10'b0011111011;
    16'b0001100000010010: out_v[177] = 10'b1101000101;
    16'b0000101010010010: out_v[177] = 10'b1001000011;
    16'b0000101100010010: out_v[177] = 10'b0110110101;
    16'b1001000000001000: out_v[177] = 10'b1000111010;
    16'b0001101100000010: out_v[177] = 10'b0100110011;
    16'b0001101100010010: out_v[177] = 10'b1110100101;
    16'b0010101010000010: out_v[177] = 10'b1000100010;
    16'b0001000100010000: out_v[177] = 10'b1010100100;
    16'b0000101110010010: out_v[177] = 10'b1110100110;
    16'b0001001100010010: out_v[177] = 10'b1010000110;
    16'b0000100010000010: out_v[177] = 10'b1000110110;
    16'b0000001010000010: out_v[177] = 10'b1101101010;
    16'b0001101100000000: out_v[177] = 10'b1010110111;
    16'b0000000100010000: out_v[177] = 10'b1011110001;
    16'b0001000100000010: out_v[177] = 10'b0111101101;
    16'b0010101000010010: out_v[177] = 10'b0011111011;
    16'b0001001100000010: out_v[177] = 10'b1001101100;
    16'b0001101000000010: out_v[177] = 10'b0101111010;
    16'b0000101110010000: out_v[177] = 10'b0110110111;
    16'b0000101100010000: out_v[177] = 10'b1011100100;
    16'b1001101100010000: out_v[177] = 10'b0011011011;
    16'b1001101110010010: out_v[177] = 10'b1111000110;
    16'b1001101110010000: out_v[177] = 10'b1011111100;
    16'b0001101100010000: out_v[177] = 10'b0101110100;
    16'b1010101010000010: out_v[177] = 10'b0011101011;
    16'b1011001010010010: out_v[177] = 10'b1111101100;
    16'b0010001010000010: out_v[177] = 10'b0110100110;
    16'b1000100110000000: out_v[177] = 10'b0111111011;
    16'b1011101110010010: out_v[177] = 10'b0111110000;
    16'b1011101010010010: out_v[177] = 10'b1011011111;
    16'b1010001010000010: out_v[177] = 10'b1010010111;
    16'b1001100110010000: out_v[177] = 10'b0011100110;
    16'b1000100110010000: out_v[177] = 10'b1011001101;
    16'b1000101110010000: out_v[177] = 10'b1011010110;
    16'b1010000010000010: out_v[177] = 10'b1110110111;
    16'b1011001010000010: out_v[177] = 10'b0110111111;
    16'b0000100100010000: out_v[177] = 10'b0110110001;
    16'b1000100010000000: out_v[177] = 10'b1011101101;
    16'b1000001010000010: out_v[177] = 10'b1000111100;
    16'b1000101100010000: out_v[177] = 10'b1011010101;
    16'b1001001000001000: out_v[177] = 10'b1111011110;
    16'b0001001010000010: out_v[177] = 10'b0111011011;
    16'b0011001010000010: out_v[177] = 10'b1111111011;
    16'b1011000010010010: out_v[177] = 10'b0011111111;
    16'b1001100110000000: out_v[177] = 10'b0110111000;
    16'b1011000010000010: out_v[177] = 10'b1111101101;
    16'b0011001010010010: out_v[177] = 10'b0011101000;
    16'b1001101110000000: out_v[177] = 10'b0111100101;
    16'b1010101110000010: out_v[177] = 10'b0111010110;
    16'b0001000100001010: out_v[177] = 10'b1011000011;
    16'b0001000110001010: out_v[177] = 10'b0100011111;
    16'b0001000100011010: out_v[177] = 10'b0011010011;
    16'b0000001110011010: out_v[177] = 10'b1011001101;
    16'b0001001110011010: out_v[177] = 10'b1010000100;
    16'b0000000010011010: out_v[177] = 10'b0011100011;
    16'b0000001010001010: out_v[177] = 10'b1011110110;
    16'b0001001110111010: out_v[177] = 10'b0111000110;
    16'b0001001100011010: out_v[177] = 10'b0110111111;
    16'b0001000110010010: out_v[177] = 10'b1000000110;
    16'b0001000100010010: out_v[177] = 10'b0010101110;
    16'b0001000110111010: out_v[177] = 10'b0101100001;
    16'b0000000110011010: out_v[177] = 10'b0011011010;
    16'b0001001110010010: out_v[177] = 10'b1111010110;
    16'b1001101000001010: out_v[177] = 10'b0111101001;
    16'b1001101100001010: out_v[177] = 10'b0111010100;
    16'b1001101100011010: out_v[177] = 10'b1011111100;
    16'b0001101100001010: out_v[177] = 10'b1011110011;
    16'b0001100100001000: out_v[177] = 10'b1001101101;
    16'b0001001000001010: out_v[177] = 10'b0101100000;
    16'b0001101000001010: out_v[177] = 10'b1110000111;
    16'b0001101100011010: out_v[177] = 10'b0111110000;
    16'b0001001100001010: out_v[177] = 10'b0100011010;
    16'b1001100100001010: out_v[177] = 10'b0010110101;
    16'b1001100000001010: out_v[177] = 10'b1010110110;
    16'b1000100100001000: out_v[177] = 10'b0100101101;
    16'b0001100000001010: out_v[177] = 10'b0101001111;
    16'b0001101000001000: out_v[177] = 10'b1110001111;
    16'b0000101000011010: out_v[177] = 10'b1011010111;
    16'b0001001000000010: out_v[177] = 10'b1101001111;
    16'b0001100100001010: out_v[177] = 10'b0001101011;
    16'b1001100100001000: out_v[177] = 10'b1110110000;
    16'b1001101100001000: out_v[177] = 10'b1110110110;
    16'b1000101000011010: out_v[177] = 10'b0110010011;
    16'b0000100100001000: out_v[177] = 10'b0111100000;
    16'b1010101000011010: out_v[177] = 10'b1111011001;
    16'b0001101000011010: out_v[177] = 10'b1111100011;
    16'b1000000100001000: out_v[177] = 10'b0110010001;
    16'b1001100000001000: out_v[177] = 10'b1111111010;
    16'b1001001110011010: out_v[177] = 10'b1010101001;
    16'b0000001100011010: out_v[177] = 10'b0100100011;
    16'b1001000110011010: out_v[177] = 10'b1110000100;
    16'b0000000110010010: out_v[177] = 10'b1011001010;
    16'b1000001110011010: out_v[177] = 10'b0110100111;
    default: out_v[177] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1011000011101000: out_v[178] = 10'b0000000101;
    16'b0011000001011000: out_v[178] = 10'b1001000001;
    16'b1011000010111000: out_v[178] = 10'b1010100111;
    16'b0011000001001000: out_v[178] = 10'b0010110001;
    16'b1011101000100000: out_v[178] = 10'b1111001111;
    16'b0011001000010000: out_v[178] = 10'b0011101111;
    16'b1001000001011000: out_v[178] = 10'b0010011110;
    16'b0001000000010000: out_v[178] = 10'b0101001111;
    16'b1011000011001000: out_v[178] = 10'b0110110101;
    16'b1011000001011000: out_v[178] = 10'b1111110101;
    16'b1001000011111000: out_v[178] = 10'b1111001011;
    16'b1001000011011000: out_v[178] = 10'b1110001001;
    16'b1011000010101000: out_v[178] = 10'b1101001111;
    16'b0011000000010000: out_v[178] = 10'b0011101000;
    16'b0001000001001000: out_v[178] = 10'b1111000010;
    16'b0001000001011000: out_v[178] = 10'b0110010001;
    16'b1011000000101000: out_v[178] = 10'b1001100110;
    16'b1011001010110000: out_v[178] = 10'b0110011111;
    16'b1011001010100000: out_v[178] = 10'b0111011101;
    16'b1001000010111000: out_v[178] = 10'b1111011110;
    16'b0011000001000000: out_v[178] = 10'b1001100011;
    16'b0010000001011000: out_v[178] = 10'b1111000011;
    16'b0000000001011000: out_v[178] = 10'b1100100011;
    16'b1011000000001000: out_v[178] = 10'b1011011101;
    16'b1001000010101000: out_v[178] = 10'b1111001101;
    16'b0000000000010000: out_v[178] = 10'b0000100011;
    16'b0011000000001000: out_v[178] = 10'b1001100010;
    16'b1011000001001000: out_v[178] = 10'b0011101011;
    16'b1001000000011000: out_v[178] = 10'b1111111011;
    16'b0011000010101000: out_v[178] = 10'b0011011101;
    16'b1001001010110000: out_v[178] = 10'b1011011111;
    16'b1011000011011000: out_v[178] = 10'b0110100110;
    16'b0011000000011000: out_v[178] = 10'b1111101010;
    16'b1010000011000000: out_v[178] = 10'b1100001001;
    16'b0010000001000000: out_v[178] = 10'b0010011001;
    16'b1011000010100000: out_v[178] = 10'b0000001110;
    16'b1011101010111000: out_v[178] = 10'b1111100000;
    16'b1011000011100000: out_v[178] = 10'b1110101000;
    16'b1011000011111000: out_v[178] = 10'b1101000010;
    16'b1011100010111000: out_v[178] = 10'b1011111111;
    16'b1011000010001000: out_v[178] = 10'b1000010011;
    16'b1011000011000000: out_v[178] = 10'b0011111110;
    16'b0001000000011000: out_v[178] = 10'b1000111010;
    16'b0010000000000000: out_v[178] = 10'b1010001110;
    16'b0000000010000000: out_v[178] = 10'b1110110001;
    16'b0000000000000000: out_v[178] = 10'b1000101110;
    16'b1000000010000000: out_v[178] = 10'b0110100010;
    16'b1000000000100000: out_v[178] = 10'b0010100011;
    16'b0011000000000000: out_v[178] = 10'b0010100101;
    16'b0011000001010000: out_v[178] = 10'b0101101000;
    16'b1000000000000000: out_v[178] = 10'b0110110100;
    16'b1000000010100000: out_v[178] = 10'b0000100110;
    16'b0000000000100000: out_v[178] = 10'b0010111111;
    16'b1010000000100000: out_v[178] = 10'b0000011101;
    16'b0010000001001000: out_v[178] = 10'b0000011110;
    16'b1010000010100000: out_v[178] = 10'b0001111100;
    16'b1011000000000000: out_v[178] = 10'b0100110111;
    16'b0010000000100000: out_v[178] = 10'b0111100110;
    16'b1010000011100000: out_v[178] = 10'b1011001001;
    16'b1001000000110000: out_v[178] = 10'b0101010100;
    16'b1010000001100000: out_v[178] = 10'b0010110100;
    16'b1010000001101000: out_v[178] = 10'b0011110100;
    16'b1011000000100000: out_v[178] = 10'b0010100100;
    16'b0010000001100000: out_v[178] = 10'b1011010111;
    16'b1001000001111000: out_v[178] = 10'b0100011010;
    16'b1011000001101000: out_v[178] = 10'b1011001100;
    16'b0001000001111000: out_v[178] = 10'b0010010011;
    16'b0000000001000000: out_v[178] = 10'b0011100100;
    16'b0010000001101000: out_v[178] = 10'b0111011010;
    16'b0000000001001000: out_v[178] = 10'b1011001100;
    16'b0001000000000000: out_v[178] = 10'b0110001001;
    16'b1010000000000000: out_v[178] = 10'b0100001111;
    16'b0011000000100000: out_v[178] = 10'b1100100110;
    16'b0011000001101000: out_v[178] = 10'b0010011000;
    16'b1011000001111000: out_v[178] = 10'b1111000011;
    16'b1000000001100000: out_v[178] = 10'b1011000111;
    16'b0000100001001000: out_v[178] = 10'b1100101100;
    16'b1011000001100000: out_v[178] = 10'b0111001010;
    16'b0010000010000000: out_v[178] = 10'b0010011110;
    16'b1000000001101000: out_v[178] = 10'b0011000010;
    16'b1010000010000000: out_v[178] = 10'b0101011001;
    16'b0000000010100000: out_v[178] = 10'b1100101001;
    16'b1000000011100000: out_v[178] = 10'b1000101011;
    16'b1010000011101000: out_v[178] = 10'b1111000010;
    16'b1000000010100010: out_v[178] = 10'b0111011001;
    16'b0000000011100000: out_v[178] = 10'b1011100110;
    16'b0010000011100000: out_v[178] = 10'b1110011001;
    16'b1000000011100010: out_v[178] = 10'b1000011111;
    16'b1000000011000000: out_v[178] = 10'b0001101110;
    16'b1011000011110000: out_v[178] = 10'b0010011011;
    16'b0010000010100000: out_v[178] = 10'b1111101010;
    16'b1011000001000000: out_v[178] = 10'b1001100010;
    16'b1011000010010000: out_v[178] = 10'b0001111011;
    16'b1011000010110000: out_v[178] = 10'b1111011110;
    16'b1011000010000000: out_v[178] = 10'b0011110001;
    16'b1010000001000000: out_v[178] = 10'b0010111000;
    16'b1010000010100010: out_v[178] = 10'b1101000100;
    16'b1010000011100010: out_v[178] = 10'b1011101110;
    16'b0001000001010000: out_v[178] = 10'b0000011111;
    16'b0000000011000000: out_v[178] = 10'b1000010001;
    16'b0011000011011000: out_v[178] = 10'b0111001111;
    16'b0010000011000000: out_v[178] = 10'b0000110110;
    16'b1000000001000000: out_v[178] = 10'b1011010001;
    16'b0010000011001000: out_v[178] = 10'b0001010011;
    16'b1010000001001000: out_v[178] = 10'b0110010011;
    16'b1010000011001000: out_v[178] = 10'b0110100111;
    16'b0011000011000000: out_v[178] = 10'b1001010000;
    16'b0001001001011000: out_v[178] = 10'b1100101111;
    16'b0000000011001000: out_v[178] = 10'b0110111001;
    16'b0001000011011000: out_v[178] = 10'b0101111110;
    16'b0011000011001000: out_v[178] = 10'b0111011010;
    16'b1000000011001000: out_v[178] = 10'b0111010100;
    16'b1011001001101000: out_v[178] = 10'b0110101111;
    16'b0010000000010000: out_v[178] = 10'b1101100000;
    16'b1000000010010000: out_v[178] = 10'b1001010101;
    16'b0010000001010000: out_v[178] = 10'b1100100000;
    16'b1010000001010000: out_v[178] = 10'b0000101011;
    16'b1010000011010000: out_v[178] = 10'b0001110110;
    16'b0000000001010000: out_v[178] = 10'b1110100110;
    16'b1000000010110000: out_v[178] = 10'b0010110010;
    16'b1000000011110000: out_v[178] = 10'b1010101111;
    16'b0010000011010000: out_v[178] = 10'b0100101110;
    16'b0001000001000000: out_v[178] = 10'b1000111001;
    16'b1011000011010000: out_v[178] = 10'b1101100110;
    16'b1000000011010000: out_v[178] = 10'b0111011111;
    16'b1000000011101000: out_v[178] = 10'b0010101000;
    16'b1010000011110000: out_v[178] = 10'b1010110011;
    16'b1010000010010000: out_v[178] = 10'b1101100100;
    16'b1000000000001000: out_v[178] = 10'b1101010100;
    16'b1000000000101000: out_v[178] = 10'b1001001000;
    16'b1000000001001000: out_v[178] = 10'b0011010100;
    16'b0000100000001000: out_v[178] = 10'b0011110011;
    16'b0001000000001000: out_v[178] = 10'b0101101101;
    16'b1000100001101000: out_v[178] = 10'b1011011110;
    16'b1001000001001000: out_v[178] = 10'b0111010100;
    16'b0000000000001000: out_v[178] = 10'b1101100110;
    16'b1001000001101000: out_v[178] = 10'b0010111100;
    16'b0111000000010000: out_v[178] = 10'b0011011101;
    16'b0111000000000000: out_v[178] = 10'b0010110000;
    16'b0011000010000000: out_v[178] = 10'b0001011100;
    16'b1011000010000010: out_v[178] = 10'b1101011010;
    16'b0110000000000000: out_v[178] = 10'b1101010111;
    16'b0011000010010000: out_v[178] = 10'b0110110111;
    16'b0011000010000010: out_v[178] = 10'b0101101110;
    16'b1011001010000000: out_v[178] = 10'b0111001110;
    16'b1001000010000000: out_v[178] = 10'b1100010110;
    16'b0011000011010000: out_v[178] = 10'b1100110110;
    16'b1001000010010000: out_v[178] = 10'b1101011100;
    16'b1001000011010000: out_v[178] = 10'b0100011010;
    16'b0001000010010000: out_v[178] = 10'b1111000110;
    16'b1001000011110000: out_v[178] = 10'b1111001010;
    16'b1001000010100000: out_v[178] = 10'b1110000001;
    16'b0001000011010000: out_v[178] = 10'b0000111011;
    16'b0001000010000000: out_v[178] = 10'b0100010100;
    16'b0011000011100000: out_v[178] = 10'b0111000011;
    16'b0011000010001000: out_v[178] = 10'b1000010111;
    16'b0111000001000000: out_v[178] = 10'b1100000111;
    16'b0111000001010000: out_v[178] = 10'b1011011111;
    16'b1010000000001000: out_v[178] = 10'b1100101011;
    16'b0000000001100000: out_v[178] = 10'b1000100001;
    default: out_v[178] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0101100100000100: out_v[179] = 10'b0111010011;
    16'b0100100010001100: out_v[179] = 10'b0110100111;
    16'b0100100000000100: out_v[179] = 10'b0011111010;
    16'b0000000100000000: out_v[179] = 10'b1001100000;
    16'b0100000100001100: out_v[179] = 10'b1010011101;
    16'b0100000100000100: out_v[179] = 10'b0110111001;
    16'b0100100010000000: out_v[179] = 10'b1111000011;
    16'b0000100000000000: out_v[179] = 10'b0001110111;
    16'b0101100100001100: out_v[179] = 10'b1001010101;
    16'b0000000100001100: out_v[179] = 10'b1011011010;
    16'b0100000000000000: out_v[179] = 10'b1000101011;
    16'b0101101100001100: out_v[179] = 10'b0000100111;
    16'b0100100110000100: out_v[179] = 10'b1001110111;
    16'b0100100100000000: out_v[179] = 10'b0010110101;
    16'b0100100000000000: out_v[179] = 10'b0000010011;
    16'b0101100000001100: out_v[179] = 10'b1000010101;
    16'b0100000000000100: out_v[179] = 10'b1000100111;
    16'b0101100000000000: out_v[179] = 10'b1111010001;
    16'b0101000100001100: out_v[179] = 10'b1000001011;
    16'b0100000110000000: out_v[179] = 10'b1000010001;
    16'b0100100100001100: out_v[179] = 10'b0100011001;
    16'b0100100100000100: out_v[179] = 10'b1001111100;
    16'b0100000110001100: out_v[179] = 10'b1011010110;
    16'b0100100000100000: out_v[179] = 10'b1111100110;
    16'b0101100000000100: out_v[179] = 10'b0111011011;
    16'b0001000100000100: out_v[179] = 10'b0101001001;
    16'b0100100010000100: out_v[179] = 10'b0011100110;
    16'b0000100010000000: out_v[179] = 10'b1010011001;
    16'b0100100100100100: out_v[179] = 10'b1110111110;
    16'b0100000110000100: out_v[179] = 10'b0101110001;
    16'b0100100000100100: out_v[179] = 10'b0100100111;
    16'b0101000100000100: out_v[179] = 10'b1100000100;
    16'b0100100000001100: out_v[179] = 10'b0011001011;
    16'b0100000100100100: out_v[179] = 10'b1111011001;
    16'b0101101100000100: out_v[179] = 10'b0000010011;
    16'b0101000100101100: out_v[179] = 10'b1000000110;
    16'b0101100100000000: out_v[179] = 10'b1100011011;
    16'b0100000010000000: out_v[179] = 10'b1111011111;
    16'b0101001100001100: out_v[179] = 10'b0010001011;
    16'b0100000100000000: out_v[179] = 10'b1010011010;
    16'b0100100110000000: out_v[179] = 10'b0100001100;
    16'b0000000100000100: out_v[179] = 10'b0110010101;
    16'b0000101100001100: out_v[179] = 10'b1001010011;
    16'b0100001000000000: out_v[179] = 10'b1010101001;
    16'b0000001000000000: out_v[179] = 10'b1111001111;
    16'b0000001100001100: out_v[179] = 10'b1101100110;
    16'b0100101100001000: out_v[179] = 10'b1110110001;
    16'b0100001000001000: out_v[179] = 10'b1001001110;
    16'b0000000000000000: out_v[179] = 10'b1001110111;
    16'b0100101100001100: out_v[179] = 10'b0110000110;
    16'b0100001000001100: out_v[179] = 10'b1101101100;
    16'b0100001100000000: out_v[179] = 10'b0101000100;
    16'b0000101000001100: out_v[179] = 10'b1010111001;
    16'b0100101100000000: out_v[179] = 10'b0111010010;
    16'b0100101000000000: out_v[179] = 10'b0010111101;
    16'b0100101000001000: out_v[179] = 10'b1011100011;
    16'b0100101000001100: out_v[179] = 10'b1001011000;
    16'b0100000000001000: out_v[179] = 10'b0110100100;
    16'b0100001100001100: out_v[179] = 10'b1110010010;
    16'b0000100000001100: out_v[179] = 10'b0010001011;
    16'b0100001100001000: out_v[179] = 10'b0100000101;
    16'b0101001100000100: out_v[179] = 10'b0111111101;
    16'b0100000100001000: out_v[179] = 10'b1010010001;
    16'b0100001100101100: out_v[179] = 10'b0110011100;
    16'b0001001100001100: out_v[179] = 10'b0010011011;
    16'b0000001100101100: out_v[179] = 10'b1010000111;
    16'b0001001000000100: out_v[179] = 10'b0000111011;
    16'b0100001100001110: out_v[179] = 10'b0111010100;
    16'b0100101100101100: out_v[179] = 10'b0011010101;
    16'b0101101000000100: out_v[179] = 10'b1000101110;
    16'b0100100100101100: out_v[179] = 10'b1011111010;
    16'b0000100100001100: out_v[179] = 10'b1000111110;
    16'b0000001100001110: out_v[179] = 10'b1110100110;
    16'b0000001100000000: out_v[179] = 10'b1000111111;
    16'b0101001100000000: out_v[179] = 10'b0101100010;
    16'b0001001100000000: out_v[179] = 10'b1101001001;
    16'b0100001100000100: out_v[179] = 10'b0000011111;
    16'b0000001000001100: out_v[179] = 10'b0001110111;
    16'b0001101000000100: out_v[179] = 10'b1000010110;
    16'b0001001100000010: out_v[179] = 10'b1001011111;
    16'b0101001110000000: out_v[179] = 10'b0011111110;
    16'b0001001100000100: out_v[179] = 10'b0111110110;
    16'b0001100000001100: out_v[179] = 10'b0101011111;
    16'b0100101000101100: out_v[179] = 10'b0100011001;
    16'b0100001000100000: out_v[179] = 10'b0100111001;
    16'b0100001000101100: out_v[179] = 10'b1100101000;
    16'b0100100000001000: out_v[179] = 10'b1111001100;
    16'b0101101000101100: out_v[179] = 10'b1000011010;
    16'b0100000000001100: out_v[179] = 10'b0110000010;
    16'b0101101000001100: out_v[179] = 10'b1011001011;
    16'b0100101000000100: out_v[179] = 10'b0001111010;
    16'b0100000000100000: out_v[179] = 10'b0011111101;
    16'b0101100000001000: out_v[179] = 10'b1000101110;
    16'b0100100000101100: out_v[179] = 10'b0100111111;
    16'b0101101000000000: out_v[179] = 10'b1100100110;
    16'b0100001000101000: out_v[179] = 10'b0110101011;
    16'b0001001010000000: out_v[179] = 10'b1101001101;
    16'b0101001000000000: out_v[179] = 10'b0010111101;
    16'b0001101010000000: out_v[179] = 10'b1001011000;
    16'b0001001000101100: out_v[179] = 10'b0100111011;
    16'b0000000000001100: out_v[179] = 10'b0011011100;
    16'b0001101000001100: out_v[179] = 10'b0100010001;
    16'b0000001000001000: out_v[179] = 10'b0000111101;
    16'b0000001000101100: out_v[179] = 10'b1111110001;
    16'b0000001000000100: out_v[179] = 10'b1101101001;
    16'b0101101010000000: out_v[179] = 10'b0110011100;
    16'b0001001000100000: out_v[179] = 10'b0110011101;
    16'b0001001000000000: out_v[179] = 10'b0011001011;
    16'b0001001000001100: out_v[179] = 10'b0010010010;
    16'b0001000000000000: out_v[179] = 10'b0111001111;
    16'b0001001000100100: out_v[179] = 10'b0111111110;
    16'b0000101000000100: out_v[179] = 10'b1001111111;
    16'b0000000000000100: out_v[179] = 10'b1001011110;
    16'b0101001000101100: out_v[179] = 10'b1010010100;
    16'b0101001000001100: out_v[179] = 10'b1101100110;
    16'b0100001110000100: out_v[179] = 10'b0110111011;
    16'b0000101010001100: out_v[179] = 10'b1011100111;
    16'b0000000110001100: out_v[179] = 10'b1101101000;
    16'b0100001010000100: out_v[179] = 10'b0000110111;
    16'b0101100000100000: out_v[179] = 10'b0111010011;
    16'b0100101010001100: out_v[179] = 10'b0111000011;
    16'b0100101010000100: out_v[179] = 10'b1001100110;
    16'b0100101010000000: out_v[179] = 10'b1001011011;
    16'b0100001000000100: out_v[179] = 10'b1000000110;
    16'b0100101000100000: out_v[179] = 10'b1010110001;
    16'b0000001110001100: out_v[179] = 10'b0011110011;
    16'b0000001010000100: out_v[179] = 10'b1100101111;
    16'b0000001010001100: out_v[179] = 10'b0100100111;
    16'b0001100000000000: out_v[179] = 10'b1110100001;
    16'b0000000010001100: out_v[179] = 10'b1001100111;
    16'b0000101000000000: out_v[179] = 10'b1010100100;
    16'b0110001100000010: out_v[179] = 10'b0101011101;
    16'b0100000100000010: out_v[179] = 10'b0111110000;
    16'b0101000100000010: out_v[179] = 10'b1111100010;
    16'b0111001100000010: out_v[179] = 10'b1110011001;
    16'b0001000100000000: out_v[179] = 10'b1101100100;
    16'b0101000100000000: out_v[179] = 10'b1101101010;
    16'b0100001100000010: out_v[179] = 10'b0001011100;
    16'b0000001100000010: out_v[179] = 10'b1011010000;
    16'b0101001100000010: out_v[179] = 10'b1011000011;
    16'b0110000100000010: out_v[179] = 10'b1001001010;
    16'b0000001100001000: out_v[179] = 10'b1100010100;
    16'b0111000100000010: out_v[179] = 10'b1001111110;
    16'b0100001000000010: out_v[179] = 10'b1110010011;
    16'b0110001100000011: out_v[179] = 10'b0011111010;
    16'b0001001100001000: out_v[179] = 10'b1001011110;
    16'b0001000000001100: out_v[179] = 10'b0010100101;
    16'b0101100010001100: out_v[179] = 10'b0101001111;
    16'b0101000000001100: out_v[179] = 10'b0100010111;
    16'b0001100010001100: out_v[179] = 10'b0011000110;
    16'b0001000000101100: out_v[179] = 10'b0101011110;
    16'b0001100000000100: out_v[179] = 10'b0010100111;
    16'b0101000000000100: out_v[179] = 10'b0101010111;
    16'b0000000000001000: out_v[179] = 10'b1101000011;
    16'b0001000000011100: out_v[179] = 10'b1111000101;
    16'b0001000000000100: out_v[179] = 10'b1001111110;
    16'b0000100000000100: out_v[179] = 10'b1110001101;
    16'b0100000000101100: out_v[179] = 10'b0011010100;
    16'b0001000000001000: out_v[179] = 10'b0011100011;
    16'b0101100010000100: out_v[179] = 10'b0111110110;
    16'b0001000000111100: out_v[179] = 10'b1011100011;
    16'b0000101100000100: out_v[179] = 10'b1110100000;
    16'b0101101110000000: out_v[179] = 10'b0001000011;
    16'b0101101100000000: out_v[179] = 10'b0110111010;
    16'b0100101110000000: out_v[179] = 10'b1010011000;
    16'b0101101110001100: out_v[179] = 10'b0100111011;
    16'b0100101100000100: out_v[179] = 10'b0111110001;
    16'b0000101100000000: out_v[179] = 10'b0110000111;
    16'b0101101110000100: out_v[179] = 10'b1101101010;
    16'b0100101110001100: out_v[179] = 10'b0101100001;
    16'b0100101110000100: out_v[179] = 10'b1010110001;
    16'b0101101100101100: out_v[179] = 10'b0001110111;
    16'b0101000000101100: out_v[179] = 10'b1001000111;
    16'b0101001000000100: out_v[179] = 10'b0101100110;
    16'b0101001000100100: out_v[179] = 10'b1101001001;
    default: out_v[179] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1000000000001100: out_v[180] = 10'b1101110110;
    16'b0100000000100100: out_v[180] = 10'b0001001011;
    16'b1100000000101000: out_v[180] = 10'b1000100001;
    16'b1100000000001000: out_v[180] = 10'b1101011001;
    16'b0000000000001100: out_v[180] = 10'b0110011000;
    16'b1101000000101100: out_v[180] = 10'b1111111111;
    16'b0100000000001100: out_v[180] = 10'b1010000101;
    16'b0000000000100100: out_v[180] = 10'b1001010010;
    16'b1000000000101000: out_v[180] = 10'b0011011011;
    16'b1000000000101100: out_v[180] = 10'b0111000101;
    16'b0000000000000000: out_v[180] = 10'b1001011110;
    16'b0100000000000100: out_v[180] = 10'b1001110111;
    16'b0100000000101100: out_v[180] = 10'b0011001100;
    16'b0000000000000100: out_v[180] = 10'b0101110011;
    16'b1100000000101100: out_v[180] = 10'b0011100101;
    16'b1000000000000100: out_v[180] = 10'b1111011001;
    16'b0100000000101000: out_v[180] = 10'b0101101010;
    16'b0000000000001000: out_v[180] = 10'b1100010010;
    16'b0100000000001000: out_v[180] = 10'b0110100011;
    16'b1101000000101000: out_v[180] = 10'b0110100111;
    16'b1101000000101101: out_v[180] = 10'b0001100110;
    16'b1001000000101000: out_v[180] = 10'b1111001010;
    16'b1000000000001000: out_v[180] = 10'b1111000011;
    16'b1000000000000000: out_v[180] = 10'b1010101001;
    16'b0100000000110100: out_v[180] = 10'b1111010001;
    16'b1100000000001100: out_v[180] = 10'b1111000111;
    16'b1101000000101001: out_v[180] = 10'b0111010000;
    16'b0100000000100000: out_v[180] = 10'b1101011110;
    16'b0000000000101100: out_v[180] = 10'b0010011110;
    16'b1001000000101001: out_v[180] = 10'b1111000010;
    16'b1001000000101100: out_v[180] = 10'b1000101111;
    16'b0001000000000101: out_v[180] = 10'b0101000110;
    16'b0000000000000001: out_v[180] = 10'b1000000100;
    16'b1001000000000100: out_v[180] = 10'b1000011101;
    16'b1000000000000001: out_v[180] = 10'b0101110100;
    16'b0001000000000001: out_v[180] = 10'b1001011111;
    16'b1001000000001101: out_v[180] = 10'b1010100111;
    16'b1001000000000000: out_v[180] = 10'b0110110101;
    16'b0000000000100000: out_v[180] = 10'b1001000011;
    16'b0100000000000000: out_v[180] = 10'b0110110111;
    16'b0001000000000000: out_v[180] = 10'b0001000110;
    16'b1001000000000001: out_v[180] = 10'b1100110011;
    16'b0000000010000001: out_v[180] = 10'b0101100111;
    16'b1000000010001001: out_v[180] = 10'b0001100111;
    16'b1000000010001000: out_v[180] = 10'b0001101000;
    16'b0001000100000101: out_v[180] = 10'b1110001110;
    16'b1000000010000000: out_v[180] = 10'b1001100111;
    16'b1001000100001000: out_v[180] = 10'b1111011101;
    16'b1001000000001001: out_v[180] = 10'b1011001100;
    16'b1000000000001001: out_v[180] = 10'b0001001101;
    16'b1001000000001000: out_v[180] = 10'b0110110111;
    16'b0001000100000000: out_v[180] = 10'b0101001111;
    16'b0000000010000000: out_v[180] = 10'b0000110100;
    16'b1001000100000000: out_v[180] = 10'b0100111111;
    16'b1000000010000001: out_v[180] = 10'b1110001101;
    16'b0000000000000101: out_v[180] = 10'b0110000100;
    16'b0001000000000100: out_v[180] = 10'b1110110101;
    16'b1001000000000101: out_v[180] = 10'b0101000111;
    16'b1000000000100100: out_v[180] = 10'b0110100100;
    16'b1000000000100000: out_v[180] = 10'b0101001111;
    16'b1001000000001100: out_v[180] = 10'b0001110101;
    16'b0001000100000001: out_v[180] = 10'b1101011101;
    16'b1000101000000100: out_v[180] = 10'b1010011101;
    16'b1000101000001100: out_v[180] = 10'b0000101001;
    16'b1000101000001000: out_v[180] = 10'b0110101101;
    16'b1100000000100100: out_v[180] = 10'b1010011111;
    16'b1000101000000000: out_v[180] = 10'b0001010111;
    16'b1000000000011000: out_v[180] = 10'b0101011001;
    16'b0000000010001000: out_v[180] = 10'b0001011111;
    16'b0000000000010000: out_v[180] = 10'b1111101110;
    16'b0000000000101000: out_v[180] = 10'b0011111010;
    16'b0000000000011000: out_v[180] = 10'b0110111111;
    16'b1000100000001000: out_v[180] = 10'b1011110101;
    16'b0000000000010100: out_v[180] = 10'b0100110000;
    16'b1000000000011100: out_v[180] = 10'b1000100010;
    16'b0000000000011100: out_v[180] = 10'b1011001011;
    16'b1000101000011100: out_v[180] = 10'b1011110011;
    16'b0000101000010100: out_v[180] = 10'b1100111111;
    16'b1000101000011000: out_v[180] = 10'b0101110111;
    16'b1100000000100000: out_v[180] = 10'b1010110111;
    16'b0000101000001100: out_v[180] = 10'b0011110011;
    16'b1000100000001100: out_v[180] = 10'b1000101011;
    16'b0000100000001100: out_v[180] = 10'b0011101001;
    16'b0000001000001100: out_v[180] = 10'b0010011001;
    16'b1000100000000000: out_v[180] = 10'b0010110011;
    16'b0000101000000100: out_v[180] = 10'b1111000100;
    16'b1000001000001000: out_v[180] = 10'b0011100010;
    16'b1000100000000100: out_v[180] = 10'b0101101101;
    16'b1100101000001100: out_v[180] = 10'b0101101001;
    16'b1000001000001100: out_v[180] = 10'b1101011110;
    16'b1000001000000000: out_v[180] = 10'b1011101000;
    16'b0000101000000000: out_v[180] = 10'b1000100011;
    16'b0000100000000000: out_v[180] = 10'b0101000100;
    16'b0000100000000100: out_v[180] = 10'b1101010110;
    16'b0000101000001000: out_v[180] = 10'b1001011100;
    16'b0000100000001000: out_v[180] = 10'b1010001111;
    16'b1000000010001100: out_v[180] = 10'b1110100110;
    16'b0000001000000100: out_v[180] = 10'b1011000100;
    default: out_v[180] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0011000000100010: out_v[181] = 10'b1001000001;
    16'b0011010000100011: out_v[181] = 10'b0110010000;
    16'b0011010000000111: out_v[181] = 10'b0011010011;
    16'b0011010000000100: out_v[181] = 10'b0011000001;
    16'b0011000000100000: out_v[181] = 10'b1010110011;
    16'b0011010000100000: out_v[181] = 10'b0100001110;
    16'b0011010000000101: out_v[181] = 10'b0001011011;
    16'b0010010000000000: out_v[181] = 10'b0001010000;
    16'b0011010000000000: out_v[181] = 10'b1011000011;
    16'b0001010000000000: out_v[181] = 10'b1001110001;
    16'b0011010000100001: out_v[181] = 10'b1101000111;
    16'b0010010000000100: out_v[181] = 10'b1110100000;
    16'b0011010000000001: out_v[181] = 10'b0010101001;
    16'b0011010000100010: out_v[181] = 10'b0110111000;
    16'b0011010000000010: out_v[181] = 10'b1010000011;
    16'b0011000000000010: out_v[181] = 10'b0011001111;
    16'b0001010000000100: out_v[181] = 10'b0001000011;
    16'b0011010000000110: out_v[181] = 10'b1100001000;
    16'b0010010000000101: out_v[181] = 10'b1000011011;
    16'b0011000000000100: out_v[181] = 10'b0010010111;
    16'b0001010000100001: out_v[181] = 10'b0101010001;
    16'b0011010000000011: out_v[181] = 10'b0010011010;
    16'b0011000000100001: out_v[181] = 10'b0110001110;
    16'b0011000000000000: out_v[181] = 10'b0011010100;
    16'b0001000000100001: out_v[181] = 10'b0011001001;
    16'b0000010000100001: out_v[181] = 10'b1111100001;
    16'b0011000000100011: out_v[181] = 10'b0010100001;
    16'b0001010000000110: out_v[181] = 10'b1000001011;
    16'b0001000000000000: out_v[181] = 10'b0101000111;
    16'b0011010000100101: out_v[181] = 10'b0011010011;
    16'b0001000000000001: out_v[181] = 10'b0001001010;
    16'b0000000000000011: out_v[181] = 10'b0110001001;
    16'b0010000000000011: out_v[181] = 10'b1101011110;
    16'b0000000000000001: out_v[181] = 10'b0011110010;
    16'b0010000000000001: out_v[181] = 10'b1010100111;
    16'b0000000000100001: out_v[181] = 10'b0000110010;
    16'b0001000000000011: out_v[181] = 10'b0101001010;
    16'b0010000000100001: out_v[181] = 10'b1101101001;
    16'b0001000000100011: out_v[181] = 10'b0111010011;
    16'b0000000000000000: out_v[181] = 10'b1011011111;
    16'b0011000000000001: out_v[181] = 10'b1100010010;
    16'b0001010000100000: out_v[181] = 10'b0110100100;
    16'b0000010000000001: out_v[181] = 10'b0000101100;
    16'b0000010000000000: out_v[181] = 10'b1000011101;
    16'b0010010000100000: out_v[181] = 10'b0010100101;
    16'b0001000000100000: out_v[181] = 10'b1100111001;
    16'b0000010000100000: out_v[181] = 10'b0000000100;
    16'b0010010000100001: out_v[181] = 10'b0000001110;
    16'b0010000000000000: out_v[181] = 10'b1011000110;
    16'b0010010000000001: out_v[181] = 10'b1010101010;
    16'b0010000000100000: out_v[181] = 10'b0101011011;
    16'b0000000000100000: out_v[181] = 10'b1000001101;
    16'b0001000000000010: out_v[181] = 10'b0101110100;
    16'b0010000000100010: out_v[181] = 10'b0000101110;
    16'b0000000000100011: out_v[181] = 10'b0001011110;
    16'b0000000000100010: out_v[181] = 10'b0001011101;
    16'b0010000000100011: out_v[181] = 10'b1110001100;
    16'b0011000000000011: out_v[181] = 10'b1100110001;
    16'b0001010000000001: out_v[181] = 10'b1000101010;
    16'b0010000000000010: out_v[181] = 10'b0010111001;
    16'b0001000000100010: out_v[181] = 10'b1101100001;
    16'b0000010000000100: out_v[181] = 10'b0001011000;
    16'b0000000000100100: out_v[181] = 10'b0100110101;
    16'b0000010000100100: out_v[181] = 10'b0011011110;
    16'b0000000000100101: out_v[181] = 10'b0110010111;
    16'b0010000000100100: out_v[181] = 10'b0101010011;
    16'b0000000000000100: out_v[181] = 10'b1001000111;
    16'b0010010000000010: out_v[181] = 10'b1010100010;
    16'b0000000000100110: out_v[181] = 10'b0101011111;
    16'b0010010000100010: out_v[181] = 10'b0111101010;
    16'b0011000000100100: out_v[181] = 10'b1100110000;
    16'b0011000000100110: out_v[181] = 10'b1101100010;
    16'b0011000000100111: out_v[181] = 10'b0101100110;
    16'b0011000000100101: out_v[181] = 10'b1000111110;
    16'b0000010000100101: out_v[181] = 10'b0011010000;
    16'b0011000000000101: out_v[181] = 10'b0010100110;
    16'b0010000000000111: out_v[181] = 10'b0111111011;
    16'b0000000000000101: out_v[181] = 10'b0110100111;
    16'b0001000000000111: out_v[181] = 10'b1100001011;
    16'b0010000000000100: out_v[181] = 10'b1010001100;
    16'b0000000000000111: out_v[181] = 10'b1101101111;
    16'b0010000000000110: out_v[181] = 10'b0111111000;
    16'b0011000000000111: out_v[181] = 10'b0011110011;
    16'b0010000000000101: out_v[181] = 10'b0110100000;
    16'b0011000000000110: out_v[181] = 10'b0010111101;
    16'b0001000000000101: out_v[181] = 10'b0010100010;
    16'b0000000000000010: out_v[181] = 10'b0110110110;
    16'b0010010000000110: out_v[181] = 10'b1100110111;
    16'b0010000000100110: out_v[181] = 10'b1000100111;
    16'b0010010000100100: out_v[181] = 10'b0010110110;
    16'b0010000000100101: out_v[181] = 10'b1100000111;
    16'b0010010000100101: out_v[181] = 10'b1001100110;
    default: out_v[181] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000010001000: out_v[182] = 10'b1101110000;
    16'b1000000010001000: out_v[182] = 10'b1101011001;
    16'b1000000000001000: out_v[182] = 10'b1001010001;
    16'b1000000000000000: out_v[182] = 10'b1011001001;
    16'b0000000000001000: out_v[182] = 10'b1010100110;
    16'b0000000000000000: out_v[182] = 10'b1000111010;
    16'b0000000010000000: out_v[182] = 10'b0110010100;
    16'b1100000000000000: out_v[182] = 10'b1011100010;
    16'b1000000010000000: out_v[182] = 10'b0110000110;
    16'b0100000000000000: out_v[182] = 10'b0111001000;
    16'b0100000010000000: out_v[182] = 10'b0010000100;
    16'b0100000000001000: out_v[182] = 10'b0011001100;
    16'b0000000000100000: out_v[182] = 10'b1010001101;
    16'b1100000000001000: out_v[182] = 10'b1010110110;
    16'b0100000010001000: out_v[182] = 10'b0101011011;
    16'b0000001000000000: out_v[182] = 10'b0011011011;
    16'b0000000000100001: out_v[182] = 10'b0001011100;
    16'b0000000010100001: out_v[182] = 10'b1110101110;
    16'b0000000010101001: out_v[182] = 10'b1110101010;
    16'b0000000000101000: out_v[182] = 10'b0110111010;
    16'b0000000000101001: out_v[182] = 10'b0111100110;
    16'b0000000010001001: out_v[182] = 10'b1111000010;
    16'b0000000010101000: out_v[182] = 10'b1101000011;
    16'b1100000010001000: out_v[182] = 10'b1001000101;
    16'b0000000000000001: out_v[182] = 10'b0011110011;
    16'b0000000010100000: out_v[182] = 10'b0111011000;
    16'b0000000000001001: out_v[182] = 10'b1010000011;
    16'b0000000010000001: out_v[182] = 10'b1010101011;
    default: out_v[182] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000001100000101: out_v[183] = 10'b0100000001;
    16'b0010000100000101: out_v[183] = 10'b0001010001;
    16'b0000001110000101: out_v[183] = 10'b0001100111;
    16'b0000000000000101: out_v[183] = 10'b0011010101;
    16'b0000000100000101: out_v[183] = 10'b1111100000;
    16'b0010000000000001: out_v[183] = 10'b1000010011;
    16'b0010001100000000: out_v[183] = 10'b0110010110;
    16'b0000001100000001: out_v[183] = 10'b1000011000;
    16'b0010001100000101: out_v[183] = 10'b0001101111;
    16'b0000001110000001: out_v[183] = 10'b0001011110;
    16'b0000001100000100: out_v[183] = 10'b1000011011;
    16'b0000001000000101: out_v[183] = 10'b1100001011;
    16'b0010001100000001: out_v[183] = 10'b1100000111;
    16'b0000000100000100: out_v[183] = 10'b1110000111;
    16'b0000001100000000: out_v[183] = 10'b0000100100;
    16'b0000000110000101: out_v[183] = 10'b0000110101;
    16'b0000001000000100: out_v[183] = 10'b0000011111;
    16'b0010001110000001: out_v[183] = 10'b0110110011;
    16'b0000000000000001: out_v[183] = 10'b0111010101;
    16'b0000001110000100: out_v[183] = 10'b0011001101;
    16'b0010001000000001: out_v[183] = 10'b0010010111;
    16'b0010000100000000: out_v[183] = 10'b0100001111;
    16'b0010000100000001: out_v[183] = 10'b0100011111;
    16'b0010000000000101: out_v[183] = 10'b0001111101;
    16'b0000001000000001: out_v[183] = 10'b1100100010;
    16'b0000000110000100: out_v[183] = 10'b1000011101;
    16'b0000000000000100: out_v[183] = 10'b1110010101;
    16'b0000000100000001: out_v[183] = 10'b0110100110;
    16'b0010001110000101: out_v[183] = 10'b0011101101;
    16'b0000000110000000: out_v[183] = 10'b0001001011;
    16'b0000000100000000: out_v[183] = 10'b1001101010;
    16'b0000000000000000: out_v[183] = 10'b1100110000;
    16'b0000001000000000: out_v[183] = 10'b0010111100;
    16'b0000000010000000: out_v[183] = 10'b1111011100;
    16'b0000001110000000: out_v[183] = 10'b0110001110;
    16'b0000001010000000: out_v[183] = 10'b0011100101;
    16'b0000001100001000: out_v[183] = 10'b1010110011;
    16'b0000000010000100: out_v[183] = 10'b1010110100;
    16'b0000001010000100: out_v[183] = 10'b0101110100;
    16'b0000001010000001: out_v[183] = 10'b0011110100;
    16'b0000000110000001: out_v[183] = 10'b0100110001;
    16'b0000001000001000: out_v[183] = 10'b0100010011;
    16'b0000001010000101: out_v[183] = 10'b0000100101;
    16'b0000000000001000: out_v[183] = 10'b1011000110;
    16'b0100000000000000: out_v[183] = 10'b0001101000;
    16'b0100001000000000: out_v[183] = 10'b0110000110;
    16'b0100000000000001: out_v[183] = 10'b0011111000;
    16'b0100001000000001: out_v[183] = 10'b1111001000;
    16'b0100000000000101: out_v[183] = 10'b0110011000;
    16'b0000000010000001: out_v[183] = 10'b1011111010;
    16'b0000000010000101: out_v[183] = 10'b0100111011;
    16'b0100001100000001: out_v[183] = 10'b0101011110;
    16'b0100000100000001: out_v[183] = 10'b0011110010;
    16'b0010000000000100: out_v[183] = 10'b0011111000;
    16'b0000000000001100: out_v[183] = 10'b1111000010;
    16'b0100000000000100: out_v[183] = 10'b1110010000;
    16'b0101000000000101: out_v[183] = 10'b1011010001;
    16'b0000000001000101: out_v[183] = 10'b1111010010;
    16'b0001000000000101: out_v[183] = 10'b1111111110;
    16'b0000100100000101: out_v[183] = 10'b1110110111;
    16'b0000000001000001: out_v[183] = 10'b1001110010;
    16'b0001000000000001: out_v[183] = 10'b0111010011;
    16'b0100001000000101: out_v[183] = 10'b1001001010;
    16'b0100001100000101: out_v[183] = 10'b0101011101;
    default: out_v[183] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000010010010000: out_v[184] = 10'b1011101001;
    16'b0010010010110000: out_v[184] = 10'b1001010001;
    16'b0010010010111000: out_v[184] = 10'b1001011011;
    16'b0010010000110000: out_v[184] = 10'b0111100111;
    16'b0000010000110000: out_v[184] = 10'b0011110000;
    16'b0000000010010000: out_v[184] = 10'b0110000011;
    16'b0000010010110000: out_v[184] = 10'b1000111011;
    16'b0000000010110000: out_v[184] = 10'b0110001101;
    16'b0010010010010000: out_v[184] = 10'b0101010101;
    16'b0000000010000000: out_v[184] = 10'b1111100001;
    16'b0010000000010000: out_v[184] = 10'b0100100001;
    16'b0000000000110000: out_v[184] = 10'b0001001010;
    16'b0000010010111000: out_v[184] = 10'b1110100010;
    16'b0000010010100000: out_v[184] = 10'b1100100011;
    16'b0010000010010000: out_v[184] = 10'b1010101101;
    16'b0000010000010000: out_v[184] = 10'b0001110001;
    16'b0010000010110000: out_v[184] = 10'b1000110101;
    16'b0000001000100000: out_v[184] = 10'b1001111010;
    16'b0010000010110100: out_v[184] = 10'b0011011101;
    16'b0000010000100000: out_v[184] = 10'b0111001001;
    16'b0010000000110000: out_v[184] = 10'b0101111101;
    16'b0100010000110000: out_v[184] = 10'b1010101000;
    16'b0010000000100000: out_v[184] = 10'b0100011001;
    16'b0010010000010000: out_v[184] = 10'b1010100000;
    16'b0000000000010000: out_v[184] = 10'b1101010100;
    16'b0010010010110100: out_v[184] = 10'b0000110010;
    16'b0010001010100000: out_v[184] = 10'b1100100111;
    16'b0010000010000000: out_v[184] = 10'b1011100010;
    16'b0010010010100000: out_v[184] = 10'b1001001001;
    16'b0000000000100000: out_v[184] = 10'b1100000101;
    16'b0010010000100000: out_v[184] = 10'b1011111111;
    16'b0000010000111000: out_v[184] = 10'b1011001011;
    16'b0010000010100000: out_v[184] = 10'b0010010011;
    16'b0100010010110000: out_v[184] = 10'b1000011111;
    16'b0000000000000000: out_v[184] = 10'b1000010101;
    16'b0000010010000000: out_v[184] = 10'b0101111100;
    16'b0000010000000000: out_v[184] = 10'b0111000110;
    16'b0010000000000000: out_v[184] = 10'b0100010000;
    16'b0100010000000000: out_v[184] = 10'b1111100110;
    16'b0010000000000100: out_v[184] = 10'b1001011100;
    16'b0000000000000100: out_v[184] = 10'b1001001011;
    16'b0100010000010000: out_v[184] = 10'b0010011011;
    16'b0100011010000000: out_v[184] = 10'b0011111111;
    16'b0100011010010000: out_v[184] = 10'b1110100111;
    16'b0100000000110000: out_v[184] = 10'b1111100101;
    16'b0100000010010000: out_v[184] = 10'b0110100101;
    16'b0000000000011000: out_v[184] = 10'b1111100100;
    16'b0100000000010000: out_v[184] = 10'b1111010111;
    16'b0000000010100000: out_v[184] = 10'b0110010110;
    16'b0100010010010000: out_v[184] = 10'b1001111011;
    16'b0000011000010000: out_v[184] = 10'b0101010010;
    16'b0100000010110000: out_v[184] = 10'b1110010100;
    16'b0000001010010000: out_v[184] = 10'b1010000110;
    16'b0000000000101000: out_v[184] = 10'b1010010010;
    16'b0100000010100000: out_v[184] = 10'b1110011010;
    16'b0000001000010000: out_v[184] = 10'b1011010011;
    16'b0100001010010000: out_v[184] = 10'b0110101001;
    16'b0110010010010000: out_v[184] = 10'b1010101011;
    16'b0100001000010000: out_v[184] = 10'b1010101101;
    16'b0010010000000000: out_v[184] = 10'b1011000100;
    16'b0110010000010000: out_v[184] = 10'b0001110111;
    16'b0110000000010000: out_v[184] = 10'b0110001010;
    16'b0010001000010000: out_v[184] = 10'b0100000010;
    16'b0100011000010000: out_v[184] = 10'b1001110011;
    16'b0010011000000000: out_v[184] = 10'b0010110100;
    16'b0000000000111000: out_v[184] = 10'b0001100111;
    16'b0100011000000000: out_v[184] = 10'b0010100101;
    16'b0000000010011000: out_v[184] = 10'b0111100010;
    16'b0110000010010000: out_v[184] = 10'b0111011011;
    16'b0100000000000000: out_v[184] = 10'b0000100100;
    16'b0000000010111000: out_v[184] = 10'b0010010011;
    16'b0000011000000000: out_v[184] = 10'b1111001001;
    16'b0000011010010000: out_v[184] = 10'b0100111111;
    16'b0010010010011000: out_v[184] = 10'b0000101110;
    16'b0110010000110000: out_v[184] = 10'b0111000110;
    16'b0010001010101000: out_v[184] = 10'b0110011011;
    16'b0000001010101000: out_v[184] = 10'b1111010010;
    16'b0010010000111000: out_v[184] = 10'b1011100110;
    16'b0110010010110000: out_v[184] = 10'b0111000101;
    16'b0010010000011000: out_v[184] = 10'b1011111110;
    16'b0000001000111000: out_v[184] = 10'b1000110010;
    16'b0000001000011000: out_v[184] = 10'b1100110011;
    16'b0000001010011000: out_v[184] = 10'b0001111001;
    16'b0000010011010000: out_v[184] = 10'b1111000001;
    16'b0000001000101000: out_v[184] = 10'b0110011010;
    16'b0000010000011000: out_v[184] = 10'b0010111111;
    16'b0000010001010000: out_v[184] = 10'b1101100010;
    16'b0000000000100100: out_v[184] = 10'b1111101010;
    16'b0010000000100100: out_v[184] = 10'b1011011001;
    16'b0000001000000000: out_v[184] = 10'b1001011111;
    16'b0000010000010100: out_v[184] = 10'b1010000111;
    16'b0000000000010100: out_v[184] = 10'b0100010111;
    16'b0010010010010100: out_v[184] = 10'b1010111011;
    16'b0010010000010100: out_v[184] = 10'b0100101001;
    16'b0010000010000100: out_v[184] = 10'b0101101001;
    16'b0000000010010100: out_v[184] = 10'b1111000110;
    16'b0010001000100000: out_v[184] = 10'b0100100001;
    16'b0000010010010100: out_v[184] = 10'b1000100110;
    16'b0010000010010100: out_v[184] = 10'b0011110101;
    16'b0010000000010100: out_v[184] = 10'b0111011010;
    16'b0100010000111000: out_v[184] = 10'b0110011011;
    16'b0100010000100000: out_v[184] = 10'b1011001010;
    16'b0010000010011000: out_v[184] = 10'b1111010001;
    16'b0000000010001000: out_v[184] = 10'b0101110101;
    16'b0000010010011000: out_v[184] = 10'b1000110010;
    16'b0000000000001000: out_v[184] = 10'b1010101010;
    16'b0000010011011000: out_v[184] = 10'b0010110010;
    16'b0010000010001000: out_v[184] = 10'b1011111010;
    16'b0000010001011000: out_v[184] = 10'b0011100011;
    16'b0000000010101000: out_v[184] = 10'b0101001001;
    16'b0010010010000000: out_v[184] = 10'b1001010111;
    16'b0000000011010000: out_v[184] = 10'b1111101000;
    16'b0000000001010000: out_v[184] = 10'b1100000011;
    default: out_v[184] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001000011110101: out_v[185] = 10'b1110000001;
    16'b0100000010110100: out_v[185] = 10'b0010110100;
    16'b0101000010100101: out_v[185] = 10'b1100011001;
    16'b0001000000000001: out_v[185] = 10'b1011011011;
    16'b0000000010110100: out_v[185] = 10'b1001110111;
    16'b0000010000110100: out_v[185] = 10'b0101110001;
    16'b0001000010100000: out_v[185] = 10'b1001110111;
    16'b0001000010110100: out_v[185] = 10'b0100110001;
    16'b0000000011110100: out_v[185] = 10'b1100010000;
    16'b0101000001110101: out_v[185] = 10'b0011010111;
    16'b0100010000110101: out_v[185] = 10'b1110110111;
    16'b0100010011110101: out_v[185] = 10'b0011111111;
    16'b0001000010100001: out_v[185] = 10'b0110111010;
    16'b0101000000110101: out_v[185] = 10'b1110100011;
    16'b0100010010110101: out_v[185] = 10'b1111001011;
    16'b0101000011110100: out_v[185] = 10'b1111011011;
    16'b0101000010110100: out_v[185] = 10'b0001110100;
    16'b0100010000010101: out_v[185] = 10'b0101001111;
    16'b0000000010110101: out_v[185] = 10'b0001001011;
    16'b0000010000110101: out_v[185] = 10'b1000100011;
    16'b0100000010110101: out_v[185] = 10'b1101101001;
    16'b0000010011110100: out_v[185] = 10'b0110011001;
    16'b0101000010110101: out_v[185] = 10'b1001010110;
    16'b0001000010110101: out_v[185] = 10'b0001111010;
    16'b0001000010100100: out_v[185] = 10'b0110001111;
    16'b0000010010110100: out_v[185] = 10'b1101111101;
    16'b0000000011110101: out_v[185] = 10'b0101111010;
    16'b0000000000110100: out_v[185] = 10'b1100100101;
    16'b0000010000010100: out_v[185] = 10'b1011100111;
    16'b0101000010100001: out_v[185] = 10'b1000010100;
    16'b0101100010110101: out_v[185] = 10'b0010001111;
    16'b0001000011110100: out_v[185] = 10'b0011100010;
    16'b0100000011110101: out_v[185] = 10'b0110110010;
    16'b0101000000110100: out_v[185] = 10'b0100100001;
    16'b0000000010100101: out_v[185] = 10'b1011110010;
    16'b0100010001110101: out_v[185] = 10'b1011110100;
    16'b0101000010100100: out_v[185] = 10'b0011001011;
    16'b0101000011110101: out_v[185] = 10'b1101100111;
    16'b0000010011110101: out_v[185] = 10'b0111011101;
    16'b0100000000000101: out_v[185] = 10'b1100011011;
    16'b0101000010100000: out_v[185] = 10'b1000101101;
    16'b0101000000010101: out_v[185] = 10'b0010110000;
    16'b0100000000110101: out_v[185] = 10'b1001110111;
    16'b0000010010110101: out_v[185] = 10'b1100001001;
    16'b0001000010100101: out_v[185] = 10'b1101011010;
    16'b0000000000000101: out_v[185] = 10'b1111100100;
    16'b0101000000000001: out_v[185] = 10'b1101101011;
    16'b0000000010100100: out_v[185] = 10'b0111100011;
    16'b0000010001110100: out_v[185] = 10'b1110110011;
    16'b0000000000110101: out_v[185] = 10'b1011101100;
    16'b0000000000000100: out_v[185] = 10'b1101110101;
    16'b0100000000010101: out_v[185] = 10'b1001010111;
    16'b0100000000110100: out_v[185] = 10'b1111001010;
    16'b0000010001110101: out_v[185] = 10'b0101001010;
    16'b0000100000110001: out_v[185] = 10'b0001000000;
    16'b0000100001110001: out_v[185] = 10'b0011111111;
    16'b0000100000000100: out_v[185] = 10'b1110110000;
    16'b0000100000010100: out_v[185] = 10'b1001000011;
    16'b0000110000000000: out_v[185] = 10'b0101001011;
    16'b0000100000010001: out_v[185] = 10'b1111100011;
    16'b0001100000000100: out_v[185] = 10'b1011000101;
    16'b0000100000100001: out_v[185] = 10'b1111010000;
    16'b0001110000000000: out_v[185] = 10'b1010000011;
    16'b0000100010100001: out_v[185] = 10'b0111111010;
    16'b0000100001010101: out_v[185] = 10'b0011110010;
    16'b0000110000000100: out_v[185] = 10'b1000000011;
    16'b0001100000000000: out_v[185] = 10'b0000011110;
    16'b0000100000010101: out_v[185] = 10'b1111011011;
    16'b0000100001100001: out_v[185] = 10'b1011110000;
    16'b0000100001110101: out_v[185] = 10'b1000010111;
    16'b0000100000000101: out_v[185] = 10'b0100111010;
    16'b0000100000110101: out_v[185] = 10'b1010100111;
    16'b0001100000010101: out_v[185] = 10'b1110000010;
    16'b0000100000010000: out_v[185] = 10'b1111100110;
    16'b0000100000000000: out_v[185] = 10'b1000001100;
    16'b0000100010000001: out_v[185] = 10'b1011100010;
    16'b0000100001010100: out_v[185] = 10'b1010010111;
    16'b0100100010100001: out_v[185] = 10'b1100010110;
    16'b0000100001010001: out_v[185] = 10'b1001100110;
    16'b0001100000010100: out_v[185] = 10'b1010101101;
    16'b0001110000000100: out_v[185] = 10'b1100101001;
    16'b0001100010100101: out_v[185] = 10'b1011100100;
    16'b0101100000000001: out_v[185] = 10'b1100000111;
    16'b0000100010100101: out_v[185] = 10'b0001101111;
    16'b0101100000100101: out_v[185] = 10'b1111100110;
    16'b0101100010100001: out_v[185] = 10'b1010011001;
    16'b0000100000000001: out_v[185] = 10'b0001100100;
    16'b0000110000010101: out_v[185] = 10'b0101100011;
    16'b0001100000110101: out_v[185] = 10'b0110011001;
    16'b0101000000000000: out_v[185] = 10'b1111101000;
    16'b0101100010000001: out_v[185] = 10'b1010110110;
    16'b0101100010100000: out_v[185] = 10'b1000101110;
    16'b0101100010100101: out_v[185] = 10'b0001001000;
    16'b0001100000000001: out_v[185] = 10'b1001100110;
    16'b0101100000000000: out_v[185] = 10'b0011011011;
    16'b0101100010110100: out_v[185] = 10'b1011111100;
    16'b0001100010100001: out_v[185] = 10'b0011011100;
    16'b0001100010000001: out_v[185] = 10'b0011110101;
    16'b0101000010000001: out_v[185] = 10'b1100111110;
    16'b0000100010110101: out_v[185] = 10'b0011011101;
    16'b0101100010000000: out_v[185] = 10'b0011001111;
    16'b0000110000110101: out_v[185] = 10'b0101000001;
    16'b0000100000100101: out_v[185] = 10'b1011101110;
    16'b0001100000100101: out_v[185] = 10'b0111001010;
    16'b0101000000100001: out_v[185] = 10'b0111000000;
    16'b0001000000100001: out_v[185] = 10'b1010011100;
    16'b0101000000100101: out_v[185] = 10'b1000000101;
    16'b0101000010000000: out_v[185] = 10'b0011101000;
    16'b0101100000110101: out_v[185] = 10'b0010011111;
    16'b0001000000110101: out_v[185] = 10'b1001001111;
    16'b0001000000000000: out_v[185] = 10'b0000010111;
    16'b0001100000100001: out_v[185] = 10'b1110101001;
    16'b0001000000100101: out_v[185] = 10'b1001011111;
    16'b0100000010100000: out_v[185] = 10'b0010010101;
    16'b0000110011110101: out_v[185] = 10'b0101100000;
    16'b0100100010110101: out_v[185] = 10'b0110001100;
    16'b0100100010110100: out_v[185] = 10'b0110011000;
    16'b0000110001010101: out_v[185] = 10'b1101010110;
    16'b0001100010110101: out_v[185] = 10'b0111000101;
    16'b0001100001110101: out_v[185] = 10'b0111001001;
    16'b0000110001110101: out_v[185] = 10'b0010000101;
    16'b0001100011110101: out_v[185] = 10'b0010111111;
    16'b0000110001010001: out_v[185] = 10'b0011101111;
    16'b0000110001110001: out_v[185] = 10'b1111000111;
    16'b0001110001010101: out_v[185] = 10'b0010011010;
    16'b0000100011110101: out_v[185] = 10'b0000011001;
    16'b0101100011110101: out_v[185] = 10'b1011111110;
    16'b0001100001010101: out_v[185] = 10'b0001011011;
    16'b0000110010110101: out_v[185] = 10'b0000011111;
    16'b0100100001110101: out_v[185] = 10'b0111001100;
    16'b0001110001110101: out_v[185] = 10'b0011110111;
    16'b0100110010110101: out_v[185] = 10'b1011011110;
    16'b0000110000010100: out_v[185] = 10'b1011000010;
    16'b0000110001010100: out_v[185] = 10'b1011001010;
    16'b0101100001110101: out_v[185] = 10'b1101100010;
    16'b0101100011110100: out_v[185] = 10'b1001100110;
    16'b0100110011110101: out_v[185] = 10'b1011011111;
    16'b0100110001110101: out_v[185] = 10'b1001011000;
    16'b0101110000000001: out_v[185] = 10'b0001011101;
    16'b0001010000000001: out_v[185] = 10'b0010011010;
    16'b0000000000000001: out_v[185] = 10'b1000111001;
    16'b0101100001010100: out_v[185] = 10'b0000010110;
    16'b0001110000000001: out_v[185] = 10'b0111110001;
    16'b0100100000000000: out_v[185] = 10'b1010011111;
    16'b0101100001110100: out_v[185] = 10'b0111111111;
    16'b0000000000010101: out_v[185] = 10'b0000010110;
    16'b0101100001010101: out_v[185] = 10'b1101000110;
    16'b0101000000010100: out_v[185] = 10'b0011001111;
    16'b0101100000010101: out_v[185] = 10'b1000010001;
    16'b0100000000000000: out_v[185] = 10'b0111011000;
    16'b0101100000010100: out_v[185] = 10'b0110111011;
    16'b0101110000000000: out_v[185] = 10'b1010000101;
    16'b0100000000000001: out_v[185] = 10'b1100010011;
    16'b0100010000000000: out_v[185] = 10'b1011011001;
    16'b0001000000010101: out_v[185] = 10'b0010011001;
    16'b0100100000100000: out_v[185] = 10'b1001111010;
    16'b0001000000000101: out_v[185] = 10'b0011100011;
    16'b0100110000000000: out_v[185] = 10'b1011011011;
    16'b0001100000000101: out_v[185] = 10'b1001110100;
    16'b0101000000000100: out_v[185] = 10'b1101111010;
    16'b0101010000000000: out_v[185] = 10'b1110101010;
    16'b0101000001010100: out_v[185] = 10'b1010010010;
    16'b0100100000000001: out_v[185] = 10'b1111001000;
    16'b0101010000000001: out_v[185] = 10'b1000000010;
    16'b0101000000000101: out_v[185] = 10'b1101101011;
    16'b0101100000000100: out_v[185] = 10'b1110001111;
    16'b0100000000100000: out_v[185] = 10'b1010011011;
    16'b0001000001010101: out_v[185] = 10'b0010011001;
    16'b0100110000000001: out_v[185] = 10'b1001011011;
    16'b0101100000000101: out_v[185] = 10'b1011100100;
    16'b0100100001010101: out_v[185] = 10'b0111110101;
    16'b0000110001110100: out_v[185] = 10'b1010110101;
    16'b0001110011110101: out_v[185] = 10'b1011110111;
    16'b0000110001010000: out_v[185] = 10'b0101110111;
    16'b0001100001110100: out_v[185] = 10'b0110110000;
    16'b0000100010110100: out_v[185] = 10'b1100010111;
    16'b0001100011110100: out_v[185] = 10'b0111011110;
    16'b0001100010110100: out_v[185] = 10'b0110110100;
    16'b0001100001010100: out_v[185] = 10'b0000101101;
    16'b0001100010100100: out_v[185] = 10'b1100110101;
    16'b0001100000110100: out_v[185] = 10'b0001110110;
    16'b0001110001110100: out_v[185] = 10'b1010110001;
    16'b0000110011110100: out_v[185] = 10'b1010000111;
    16'b0000100000110100: out_v[185] = 10'b1111011000;
    16'b0100010010110100: out_v[185] = 10'b1010100110;
    16'b0000110000110100: out_v[185] = 10'b1011110110;
    16'b0000100001110100: out_v[185] = 10'b1111011010;
    16'b0000110010110100: out_v[185] = 10'b1001100111;
    16'b0000110001110000: out_v[185] = 10'b0011110010;
    16'b0001000000100100: out_v[185] = 10'b0100101010;
    16'b0001000000000100: out_v[185] = 10'b1111010010;
    16'b0001000000001000: out_v[185] = 10'b0101001011;
    16'b0000000000000000: out_v[185] = 10'b0011100110;
    16'b0100100000001000: out_v[185] = 10'b1110110111;
    16'b0100000000000100: out_v[185] = 10'b1011100011;
    16'b0100000000001000: out_v[185] = 10'b1100110111;
    16'b0100100000000100: out_v[185] = 10'b1111011010;
    16'b0101000000001000: out_v[185] = 10'b0111101101;
    16'b0101100000001000: out_v[185] = 10'b0111101001;
    16'b0101100000100100: out_v[185] = 10'b1001111000;
    16'b0100100000100100: out_v[185] = 10'b1101011010;
    16'b0000100000100100: out_v[185] = 10'b0000011110;
    16'b0001100000100100: out_v[185] = 10'b1110110011;
    16'b0000000001010101: out_v[185] = 10'b0111100100;
    16'b0100010000000001: out_v[185] = 10'b0011001010;
    16'b0101000001010101: out_v[185] = 10'b1010000000;
    16'b0000000001010001: out_v[185] = 10'b0111010001;
    16'b0100000001110001: out_v[185] = 10'b0111001001;
    16'b0101010000010101: out_v[185] = 10'b0111100111;
    16'b0101000001110001: out_v[185] = 10'b0111010011;
    16'b0100000000100001: out_v[185] = 10'b0111001000;
    16'b0101010000000101: out_v[185] = 10'b0111110101;
    16'b0100000001010101: out_v[185] = 10'b0011101011;
    16'b0100000001100001: out_v[185] = 10'b0111011110;
    16'b0100000001110101: out_v[185] = 10'b1011101111;
    16'b0101000001100001: out_v[185] = 10'b0111101011;
    16'b0101110000010100: out_v[185] = 10'b0110011111;
    16'b0101110001110101: out_v[185] = 10'b1001011001;
    16'b0101110011110101: out_v[185] = 10'b1111110010;
    16'b0001110000010101: out_v[185] = 10'b0111100011;
    16'b0100100001110100: out_v[185] = 10'b0101011010;
    16'b0101110000010101: out_v[185] = 10'b0101100101;
    16'b0001110000000101: out_v[185] = 10'b0110011000;
    16'b0100100011110101: out_v[185] = 10'b1101101110;
    16'b0101100000110100: out_v[185] = 10'b1110000111;
    16'b0000110000000101: out_v[185] = 10'b0101011100;
    16'b0101110001010101: out_v[185] = 10'b1001011001;
    16'b0100100011110100: out_v[185] = 10'b0011111100;
    16'b0100110000010101: out_v[185] = 10'b0100001101;
    16'b0101110001110100: out_v[185] = 10'b0011001011;
    16'b0100110000010100: out_v[185] = 10'b0110100010;
    16'b0100100000110100: out_v[185] = 10'b1100001000;
    16'b0100110000110100: out_v[185] = 10'b1110010110;
    16'b0100100001010100: out_v[185] = 10'b1000101011;
    16'b0100100000100001: out_v[185] = 10'b1001000011;
    default: out_v[185] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100100001000000: out_v[186] = 10'b1011100000;
    16'b0100100001100000: out_v[186] = 10'b0011100111;
    16'b0100100001100010: out_v[186] = 10'b0010011011;
    16'b0000100001100010: out_v[186] = 10'b0011010110;
    16'b0000100001000000: out_v[186] = 10'b0101001001;
    16'b0001100001100010: out_v[186] = 10'b0100111100;
    16'b0001100001000000: out_v[186] = 10'b1100111011;
    16'b0100100000000000: out_v[186] = 10'b0011100001;
    16'b0000100001100000: out_v[186] = 10'b0110101011;
    16'b0000100001000010: out_v[186] = 10'b1111001111;
    16'b0001000001000010: out_v[186] = 10'b1000011001;
    16'b0000100000100000: out_v[186] = 10'b0011111010;
    16'b0001100001100000: out_v[186] = 10'b0110111111;
    16'b0001000001100010: out_v[186] = 10'b0001110111;
    16'b0000000001000010: out_v[186] = 10'b0111110011;
    16'b0000000001000000: out_v[186] = 10'b0000110111;
    16'b0100000001100000: out_v[186] = 10'b0010101001;
    16'b0001100001000010: out_v[186] = 10'b1010101111;
    16'b0101100001100010: out_v[186] = 10'b0110100111;
    16'b0001000001000000: out_v[186] = 10'b1111010001;
    16'b0101100001000000: out_v[186] = 10'b1111001101;
    16'b0000100000000000: out_v[186] = 10'b0010110001;
    16'b0001000000000010: out_v[186] = 10'b0111100111;
    16'b0001100000000000: out_v[186] = 10'b1100011011;
    16'b0101100001100000: out_v[186] = 10'b0011101010;
    16'b0100100000100000: out_v[186] = 10'b0010001010;
    16'b0100100001100100: out_v[186] = 10'b0101110110;
    16'b0101100001000010: out_v[186] = 10'b0011110110;
    16'b0100000001000100: out_v[186] = 10'b0110011010;
    16'b0000000001000100: out_v[186] = 10'b0010101110;
    16'b0000000000100100: out_v[186] = 10'b1011001100;
    16'b0100000000000100: out_v[186] = 10'b0100011000;
    16'b0100000000100100: out_v[186] = 10'b0111000011;
    16'b0100100000100100: out_v[186] = 10'b1011001101;
    16'b0000000000000100: out_v[186] = 10'b1000101110;
    16'b0100000001100100: out_v[186] = 10'b1101011010;
    16'b0000000001100100: out_v[186] = 10'b0010011110;
    16'b0000000001100000: out_v[186] = 10'b0010100110;
    16'b0001000001100000: out_v[186] = 10'b1100011111;
    16'b0000000000100000: out_v[186] = 10'b1110000100;
    16'b0000000001100101: out_v[186] = 10'b0111100101;
    16'b0000001001100100: out_v[186] = 10'b1010010110;
    16'b0000001001100000: out_v[186] = 10'b0010000110;
    16'b0000000011100100: out_v[186] = 10'b1101001000;
    16'b0000001001000100: out_v[186] = 10'b0001001110;
    16'b0000000000000000: out_v[186] = 10'b1000100000;
    16'b0000100001100100: out_v[186] = 10'b1100100010;
    16'b0001000011100100: out_v[186] = 10'b0110011011;
    16'b0001000001100100: out_v[186] = 10'b1001110110;
    16'b0001000000000100: out_v[186] = 10'b0001001111;
    16'b0001000000100100: out_v[186] = 10'b0110000110;
    16'b0100001000000100: out_v[186] = 10'b1100100111;
    16'b0100100001000100: out_v[186] = 10'b0111001010;
    16'b0100000001000000: out_v[186] = 10'b1101011000;
    16'b0100100000000100: out_v[186] = 10'b1110001101;
    16'b0100101001000100: out_v[186] = 10'b0111001000;
    16'b0000001000000100: out_v[186] = 10'b1101011011;
    16'b0100101001000000: out_v[186] = 10'b1111011010;
    16'b0100001001000100: out_v[186] = 10'b1101101011;
    16'b0100000000000000: out_v[186] = 10'b0010011011;
    16'b0000100000000100: out_v[186] = 10'b0100110000;
    16'b0100000000100000: out_v[186] = 10'b1011011001;
    16'b0000100000100100: out_v[186] = 10'b1001010001;
    16'b0000000000100110: out_v[186] = 10'b1101000100;
    16'b0000100001000100: out_v[186] = 10'b1001110010;
    16'b0000000000000010: out_v[186] = 10'b1001011011;
    16'b0000100000000110: out_v[186] = 10'b0010011101;
    16'b0000100000100110: out_v[186] = 10'b0100110111;
    16'b0000000000000110: out_v[186] = 10'b1000110001;
    16'b0000000000100010: out_v[186] = 10'b1001110011;
    16'b0000001000000110: out_v[186] = 10'b0000111010;
    16'b0100100001101000: out_v[186] = 10'b1011111110;
    16'b0100100001101100: out_v[186] = 10'b0010101110;
    16'b0100000001101100: out_v[186] = 10'b1011111000;
    16'b0000100001101100: out_v[186] = 10'b0110110010;
    16'b0000000001000110: out_v[186] = 10'b1100110000;
    16'b0001000000100110: out_v[186] = 10'b0111111000;
    16'b0001100000100000: out_v[186] = 10'b1101010010;
    16'b0101100001100100: out_v[186] = 10'b1110001101;
    16'b0001100001100100: out_v[186] = 10'b1010100001;
    16'b0001100001000100: out_v[186] = 10'b1001010010;
    16'b0001000001100110: out_v[186] = 10'b1101011010;
    16'b0001100000100100: out_v[186] = 10'b1101010011;
    16'b0100100000000010: out_v[186] = 10'b0011100100;
    16'b0100100000100010: out_v[186] = 10'b1000100110;
    16'b0000100000100010: out_v[186] = 10'b0111011000;
    16'b0000100001100110: out_v[186] = 10'b1111000010;
    16'b0100100000000110: out_v[186] = 10'b1011100110;
    default: out_v[186] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001100100010000: out_v[187] = 10'b0101010101;
    16'b0000100000010110: out_v[187] = 10'b0000111101;
    16'b0010000110010110: out_v[187] = 10'b1111110000;
    16'b0001000100010000: out_v[187] = 10'b1011001011;
    16'b0000000000010000: out_v[187] = 10'b1001101011;
    16'b0010000010010100: out_v[187] = 10'b0111011010;
    16'b0000000000010100: out_v[187] = 10'b1101110001;
    16'b0000000100010110: out_v[187] = 10'b1010110010;
    16'b0010000000010100: out_v[187] = 10'b0010001101;
    16'b0010001110010100: out_v[187] = 10'b1110110001;
    16'b0000000000010110: out_v[187] = 10'b1101000101;
    16'b0001000000010100: out_v[187] = 10'b0010110101;
    16'b0000000010010110: out_v[187] = 10'b1011010101;
    16'b0010000110010100: out_v[187] = 10'b1101010011;
    16'b0000000100010100: out_v[187] = 10'b1101011100;
    16'b0000100000000110: out_v[187] = 10'b1111000111;
    16'b0001000100010010: out_v[187] = 10'b1100010110;
    16'b0001000110010000: out_v[187] = 10'b0011101110;
    16'b0010000100010100: out_v[187] = 10'b0011100011;
    16'b0000000110010100: out_v[187] = 10'b1110001111;
    16'b0001000000010110: out_v[187] = 10'b1000101000;
    16'b0000000000010010: out_v[187] = 10'b1000100101;
    16'b0011001110010000: out_v[187] = 10'b1100100101;
    16'b0011001110010100: out_v[187] = 10'b0100000110;
    16'b0010101110010100: out_v[187] = 10'b0110011011;
    16'b0000000010010100: out_v[187] = 10'b1011101111;
    16'b0010101110000100: out_v[187] = 10'b1101000011;
    16'b0010001110010110: out_v[187] = 10'b1110100111;
    16'b0001000000010000: out_v[187] = 10'b1101001011;
    16'b0000100100000000: out_v[187] = 10'b0010011100;
    16'b0010000100010110: out_v[187] = 10'b1101110011;
    16'b0000000100010000: out_v[187] = 10'b1010111010;
    16'b0001000000010010: out_v[187] = 10'b0111000101;
    16'b0011101110010000: out_v[187] = 10'b1110000000;
    16'b0010100110010100: out_v[187] = 10'b1001001101;
    16'b0011000110010100: out_v[187] = 10'b0011110111;
    16'b0000000110010000: out_v[187] = 10'b0001111010;
    16'b0010001100010100: out_v[187] = 10'b1101010110;
    16'b0010001110010000: out_v[187] = 10'b1010111101;
    16'b0011000110010000: out_v[187] = 10'b0010010111;
    16'b0001000100010110: out_v[187] = 10'b1010111011;
    16'b0000000000000000: out_v[187] = 10'b1100010100;
    16'b0000000100000000: out_v[187] = 10'b0111010011;
    16'b0000100000010000: out_v[187] = 10'b0111111101;
    16'b0001100000010000: out_v[187] = 10'b1101001001;
    16'b0000100000000000: out_v[187] = 10'b0001100111;
    16'b0001000000000010: out_v[187] = 10'b1101000010;
    16'b0001000000000000: out_v[187] = 10'b1000001111;
    16'b0101000110010000: out_v[187] = 10'b1110010011;
    16'b0001001110010000: out_v[187] = 10'b0110100110;
    16'b0001010000010000: out_v[187] = 10'b1010101100;
    16'b0001000010010110: out_v[187] = 10'b1011010010;
    16'b0001010110010000: out_v[187] = 10'b1011000101;
    16'b0001000000000110: out_v[187] = 10'b1010100101;
    16'b0001000000000100: out_v[187] = 10'b0000101111;
    16'b0010001100010000: out_v[187] = 10'b1011110111;
    16'b0001000110010110: out_v[187] = 10'b1101100111;
    16'b0000010000010100: out_v[187] = 10'b0101001001;
    16'b0001000110000110: out_v[187] = 10'b0110101111;
    16'b0001000010000110: out_v[187] = 10'b0110111000;
    16'b0001000110000100: out_v[187] = 10'b1011111111;
    16'b0011001100010000: out_v[187] = 10'b0000101111;
    16'b0000001100010100: out_v[187] = 10'b1000001010;
    16'b0001000100000110: out_v[187] = 10'b0110110111;
    16'b0001000110010010: out_v[187] = 10'b0111011010;
    16'b0011000000000000: out_v[187] = 10'b0011100111;
    16'b0000000110010110: out_v[187] = 10'b1110100111;
    16'b0011001110010010: out_v[187] = 10'b1111010100;
    16'b0001000100000100: out_v[187] = 10'b0111011010;
    16'b0001001100000000: out_v[187] = 10'b0100101110;
    16'b0001000100010100: out_v[187] = 10'b1111100010;
    16'b0000001110010000: out_v[187] = 10'b1010001010;
    16'b0001010010010000: out_v[187] = 10'b0110011101;
    16'b0001000010010000: out_v[187] = 10'b0011000111;
    16'b0001000110010100: out_v[187] = 10'b1110100001;
    16'b0001001110010100: out_v[187] = 10'b1011111110;
    16'b0000001100010000: out_v[187] = 10'b1100010011;
    16'b0001001100010000: out_v[187] = 10'b1101111110;
    16'b0001010110010100: out_v[187] = 10'b1100110111;
    16'b0001010100010000: out_v[187] = 10'b0111000010;
    16'b0011001110010110: out_v[187] = 10'b0010001111;
    16'b0001000100000000: out_v[187] = 10'b0001110110;
    16'b0010101100000000: out_v[187] = 10'b1100001011;
    16'b0000000100010010: out_v[187] = 10'b1100100010;
    16'b0000100110000000: out_v[187] = 10'b1010001100;
    16'b0000101110010000: out_v[187] = 10'b0000011110;
    16'b0010101110000000: out_v[187] = 10'b0011111110;
    16'b0000001100000000: out_v[187] = 10'b1110101111;
    16'b0000101100000000: out_v[187] = 10'b0011001011;
    16'b0000101110000000: out_v[187] = 10'b1001100100;
    16'b0010101100010000: out_v[187] = 10'b0011111100;
    16'b0000100100010000: out_v[187] = 10'b1110100010;
    16'b0000001100010010: out_v[187] = 10'b1110010100;
    16'b0000100100010010: out_v[187] = 10'b1011010110;
    16'b0010101110010000: out_v[187] = 10'b1001111100;
    16'b0000101100010000: out_v[187] = 10'b0101101110;
    16'b0000001110000000: out_v[187] = 10'b1101100001;
    16'b0000000010010000: out_v[187] = 10'b0001101111;
    16'b0010001110000000: out_v[187] = 10'b0110000001;
    16'b0010100100000000: out_v[187] = 10'b1001011111;
    16'b0000000110000000: out_v[187] = 10'b1101101010;
    16'b0000001110010100: out_v[187] = 10'b1001101010;
    16'b0000100100000010: out_v[187] = 10'b1011001100;
    16'b0000010000010000: out_v[187] = 10'b1100011001;
    16'b0011001000000000: out_v[187] = 10'b0011111011;
    16'b0010000000000000: out_v[187] = 10'b0011011000;
    16'b0010001000000000: out_v[187] = 10'b0010110110;
    16'b0000100000010010: out_v[187] = 10'b0110111001;
    16'b0010001010000000: out_v[187] = 10'b1001010111;
    16'b0000000000000010: out_v[187] = 10'b1101100101;
    16'b0000000100000010: out_v[187] = 10'b0110101000;
    16'b0010000100000000: out_v[187] = 10'b0011000011;
    16'b0010001100000000: out_v[187] = 10'b1101100001;
    16'b0000100000000010: out_v[187] = 10'b0000101010;
    16'b0010001000000010: out_v[187] = 10'b1111000110;
    16'b0010100000010000: out_v[187] = 10'b0111011001;
    16'b0000000010000000: out_v[187] = 10'b0011011010;
    16'b0010000000000010: out_v[187] = 10'b0011110110;
    16'b0010000010000000: out_v[187] = 10'b0100010100;
    16'b0000001000000000: out_v[187] = 10'b0011010001;
    16'b0000000000000100: out_v[187] = 10'b0101011001;
    16'b0010100000000000: out_v[187] = 10'b0010011010;
    16'b0010101110010010: out_v[187] = 10'b0111010111;
    16'b0000100110000010: out_v[187] = 10'b1010101011;
    16'b0010000110010010: out_v[187] = 10'b1101100111;
    16'b0010101100010010: out_v[187] = 10'b1111101011;
    16'b0000000110010010: out_v[187] = 10'b0011110110;
    16'b0010001110010010: out_v[187] = 10'b1011111110;
    16'b0010000000010000: out_v[187] = 10'b1110111010;
    16'b0000010100010000: out_v[187] = 10'b1011100011;
    16'b0011010100010000: out_v[187] = 10'b1010011001;
    16'b0011001010010000: out_v[187] = 10'b0100000111;
    16'b0001010100000000: out_v[187] = 10'b1110101101;
    16'b0011010110010000: out_v[187] = 10'b1111011110;
    16'b0000010100000000: out_v[187] = 10'b1111000110;
    16'b0011001000010000: out_v[187] = 10'b0011011011;
    16'b0001010110000000: out_v[187] = 10'b1110010111;
    16'b0001000010010010: out_v[187] = 10'b0101000000;
    16'b0011011110010000: out_v[187] = 10'b1010001011;
    16'b0011001010000000: out_v[187] = 10'b0010010001;
    16'b0010000000000001: out_v[187] = 10'b1110011001;
    16'b0010101000000000: out_v[187] = 10'b0011110100;
    16'b0010101000010000: out_v[187] = 10'b1110100011;
    16'b0000101000010000: out_v[187] = 10'b0111000001;
    16'b0000101000000000: out_v[187] = 10'b1110010001;
    16'b0010001000010000: out_v[187] = 10'b1101111101;
    16'b0011101100000000: out_v[187] = 10'b0111111010;
    16'b0001100000000000: out_v[187] = 10'b1100000000;
    16'b0001100000010010: out_v[187] = 10'b0011000010;
    16'b0001100000000010: out_v[187] = 10'b1110000111;
    16'b0001100100000010: out_v[187] = 10'b1010110011;
    16'b0001100100010010: out_v[187] = 10'b1010001011;
    16'b0011100100010000: out_v[187] = 10'b0101000101;
    16'b0010100100010000: out_v[187] = 10'b1101001010;
    16'b0011101100010000: out_v[187] = 10'b0101000110;
    16'b0011101100010010: out_v[187] = 10'b0001010010;
    16'b0011100000010000: out_v[187] = 10'b0111000010;
    16'b0011000100010000: out_v[187] = 10'b1011101100;
    16'b0011100100010010: out_v[187] = 10'b1011110101;
    16'b0001100100000000: out_v[187] = 10'b0100110011;
    16'b0011100100000010: out_v[187] = 10'b0101110011;
    16'b0011000100000000: out_v[187] = 10'b1001101011;
    16'b0011000000000100: out_v[187] = 10'b1000100111;
    16'b0011001100000000: out_v[187] = 10'b1001101011;
    16'b0011001110000000: out_v[187] = 10'b1011000011;
    default: out_v[187] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000000010000: out_v[188] = 10'b0011110011;
    16'b1000000001010000: out_v[188] = 10'b0110111001;
    16'b0000010000010000: out_v[188] = 10'b1010100001;
    16'b0100001100001000: out_v[188] = 10'b0011111001;
    16'b0000000100010110: out_v[188] = 10'b1011001001;
    16'b0100001000001000: out_v[188] = 10'b0001101010;
    16'b1100011100001000: out_v[188] = 10'b0111100010;
    16'b0100011100001000: out_v[188] = 10'b0001101011;
    16'b1000000000010000: out_v[188] = 10'b1110101000;
    16'b1100001100001000: out_v[188] = 10'b1011110100;
    16'b1000010000010000: out_v[188] = 10'b0101101001;
    16'b0100001100000000: out_v[188] = 10'b1100100001;
    16'b0000010100010000: out_v[188] = 10'b0111010011;
    16'b1000000101010000: out_v[188] = 10'b0110111001;
    16'b0100011100000000: out_v[188] = 10'b0110000111;
    16'b1100001100011000: out_v[188] = 10'b1111011001;
    16'b1000000000000000: out_v[188] = 10'b1110110111;
    16'b0100001100011000: out_v[188] = 10'b0011111101;
    16'b0000000100010000: out_v[188] = 10'b1010100010;
    16'b1000010100010000: out_v[188] = 10'b0111100011;
    16'b0000010100000000: out_v[188] = 10'b0101001110;
    16'b0100000100011000: out_v[188] = 10'b1010001001;
    16'b0100001100001110: out_v[188] = 10'b0101010101;
    16'b0000000000000000: out_v[188] = 10'b0110000000;
    16'b1100001100001110: out_v[188] = 10'b0101110001;
    16'b1100001101001000: out_v[188] = 10'b1110010001;
    16'b1000000100010000: out_v[188] = 10'b0101110100;
    16'b1000000100010110: out_v[188] = 10'b0001011011;
    16'b0100001100011110: out_v[188] = 10'b0010111010;
    16'b0000010000000000: out_v[188] = 10'b1101000011;
    16'b0100010100000000: out_v[188] = 10'b1111111010;
    16'b0100001100010000: out_v[188] = 10'b0010111001;
    16'b0100011100010000: out_v[188] = 10'b0111101011;
    16'b0000000100000000: out_v[188] = 10'b0100010000;
    16'b0000000001000000: out_v[188] = 10'b0000011111;
    16'b1000000001000000: out_v[188] = 10'b0100001011;
    16'b0100011000010000: out_v[188] = 10'b0111011100;
    16'b1000010000000000: out_v[188] = 10'b0001011110;
    16'b1100011000000000: out_v[188] = 10'b1011011011;
    16'b0000011000000000: out_v[188] = 10'b1000100110;
    16'b0100001000000000: out_v[188] = 10'b0000011011;
    16'b0100001000010000: out_v[188] = 10'b1100001101;
    16'b0000010000000110: out_v[188] = 10'b1010001011;
    16'b0100011000000000: out_v[188] = 10'b0111011110;
    16'b1000010100000000: out_v[188] = 10'b0010011100;
    16'b0000001000000000: out_v[188] = 10'b0000010100;
    16'b0000011000010000: out_v[188] = 10'b1010110100;
    16'b0010000000000000: out_v[188] = 10'b0011111111;
    16'b0100000000010000: out_v[188] = 10'b1110100001;
    16'b1000011000000000: out_v[188] = 10'b1111100110;
    16'b0010010000000000: out_v[188] = 10'b1001110100;
    16'b1100011000010000: out_v[188] = 10'b0000010100;
    16'b1010010000010000: out_v[188] = 10'b1101110011;
    16'b1010010000000000: out_v[188] = 10'b1110101010;
    16'b1100001000000000: out_v[188] = 10'b0111010011;
    16'b1100001001000000: out_v[188] = 10'b1011011110;
    16'b1010000000000000: out_v[188] = 10'b1001011000;
    16'b1010000000010000: out_v[188] = 10'b1111011111;
    16'b1010000001010000: out_v[188] = 10'b1111110011;
    16'b1100001001010000: out_v[188] = 10'b1010011111;
    16'b1100001000010000: out_v[188] = 10'b0111101110;
    16'b0100000100010000: out_v[188] = 10'b0110011110;
    16'b1000000101000000: out_v[188] = 10'b1111100001;
    16'b0000000100001000: out_v[188] = 10'b0010010111;
    16'b0000000100011000: out_v[188] = 10'b0101010110;
    16'b0000000000001000: out_v[188] = 10'b0110000111;
    16'b0000000000011000: out_v[188] = 10'b1100100101;
    16'b0000000100010010: out_v[188] = 10'b1101101010;
    16'b1000000100000000: out_v[188] = 10'b1010110110;
    16'b1100001101000000: out_v[188] = 10'b1011100111;
    16'b1100001100010000: out_v[188] = 10'b0101100110;
    16'b1100001100000000: out_v[188] = 10'b1111010000;
    16'b0000100000010000: out_v[188] = 10'b0111100000;
    16'b0100000100000000: out_v[188] = 10'b1100001111;
    16'b0100010100010000: out_v[188] = 10'b1010100111;
    16'b0100011000001000: out_v[188] = 10'b0011010011;
    16'b0100010000010000: out_v[188] = 10'b1101011110;
    16'b0100011100011000: out_v[188] = 10'b1001011000;
    16'b0000100000000000: out_v[188] = 10'b1111010111;
    16'b0100010000000000: out_v[188] = 10'b1110111110;
    16'b0100010100001000: out_v[188] = 10'b0011111101;
    16'b0100000100001000: out_v[188] = 10'b1011000111;
    16'b0100000000000000: out_v[188] = 10'b1101100110;
    16'b0000000101000000: out_v[188] = 10'b1100000010;
    default: out_v[188] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000000000000: out_v[189] = 10'b0110001011;
    16'b0100000000010000: out_v[189] = 10'b0010110000;
    16'b0101000000000000: out_v[189] = 10'b0110010101;
    16'b0100000000000000: out_v[189] = 10'b0011110001;
    16'b0100000000000010: out_v[189] = 10'b1001001100;
    16'b0000000100000000: out_v[189] = 10'b0000111000;
    16'b0101000000010000: out_v[189] = 10'b0111100101;
    16'b0100000000010010: out_v[189] = 10'b1000101101;
    16'b0000000000010000: out_v[189] = 10'b0111110011;
    16'b0100000100000010: out_v[189] = 10'b0101010001;
    16'b0100000100000000: out_v[189] = 10'b1000100010;
    16'b0101000000000010: out_v[189] = 10'b0111010001;
    16'b0000000000000010: out_v[189] = 10'b1000111110;
    16'b0000000100000010: out_v[189] = 10'b0011000000;
    16'b0001000000000000: out_v[189] = 10'b0110111110;
    16'b0101000000010010: out_v[189] = 10'b1100011010;
    16'b0100000100010010: out_v[189] = 10'b0101010101;
    16'b0000001100000010: out_v[189] = 10'b1110001101;
    16'b0000000101000010: out_v[189] = 10'b1011100101;
    16'b0001000000000010: out_v[189] = 10'b1000101110;
    16'b0001000100000010: out_v[189] = 10'b0011000100;
    16'b0001000100000000: out_v[189] = 10'b1000101101;
    16'b0000010100000010: out_v[189] = 10'b1111010101;
    16'b0000001100000000: out_v[189] = 10'b1000000111;
    16'b0100001100000010: out_v[189] = 10'b1000110110;
    16'b0100000100010000: out_v[189] = 10'b1110101000;
    16'b0101000100000000: out_v[189] = 10'b1001001010;
    16'b0101000100010000: out_v[189] = 10'b1000111010;
    16'b0000000100010000: out_v[189] = 10'b1100010010;
    16'b0000000010000000: out_v[189] = 10'b0110001101;
    16'b0100000110000000: out_v[189] = 10'b0011110010;
    16'b0000000110000010: out_v[189] = 10'b1010110010;
    16'b0000000010000010: out_v[189] = 10'b0010101101;
    16'b0000000110000000: out_v[189] = 10'b0110100110;
    16'b0100010100000010: out_v[189] = 10'b0101110010;
    16'b0100010000000000: out_v[189] = 10'b1001100010;
    16'b0100010000000010: out_v[189] = 10'b0101001011;
    16'b0100000110000010: out_v[189] = 10'b1100101010;
    default: out_v[189] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000100100001000: out_v[190] = 10'b0010110001;
    16'b0000001000000010: out_v[190] = 10'b0000101110;
    16'b0000100000000010: out_v[190] = 10'b1110110001;
    16'b0000000100000000: out_v[190] = 10'b0100110100;
    16'b1000001000000110: out_v[190] = 10'b0001000000;
    16'b1000101000000110: out_v[190] = 10'b0001101010;
    16'b0000101100000000: out_v[190] = 10'b1011011000;
    16'b1000001000001110: out_v[190] = 10'b1101100011;
    16'b0000001100000000: out_v[190] = 10'b1000001011;
    16'b0000101100000010: out_v[190] = 10'b1110000100;
    16'b0000101000001010: out_v[190] = 10'b1100000111;
    16'b0000001000001010: out_v[190] = 10'b1010001001;
    16'b0000000000000000: out_v[190] = 10'b0000111111;
    16'b0000000100001000: out_v[190] = 10'b0011011000;
    16'b0000100100000000: out_v[190] = 10'b0001111001;
    16'b1000001000000010: out_v[190] = 10'b0011110100;
    16'b0000101100001010: out_v[190] = 10'b1110010011;
    16'b0000101000000010: out_v[190] = 10'b1011111000;
    16'b0000001100001000: out_v[190] = 10'b0011111100;
    16'b1000101100000110: out_v[190] = 10'b0110101001;
    16'b0000001100000010: out_v[190] = 10'b0000100011;
    16'b0000001100001010: out_v[190] = 10'b0101111000;
    16'b0000000000000010: out_v[190] = 10'b0010001011;
    16'b0000100000001010: out_v[190] = 10'b1111000110;
    16'b1000101000001110: out_v[190] = 10'b0010000001;
    16'b0000100000000000: out_v[190] = 10'b0100101101;
    16'b0000001000000000: out_v[190] = 10'b1000110100;
    16'b0000100100000010: out_v[190] = 10'b0110110101;
    16'b0000100100001010: out_v[190] = 10'b1110000011;
    16'b1000101100001110: out_v[190] = 10'b1001101011;
    16'b0000000000001010: out_v[190] = 10'b0011001011;
    16'b0000001000000110: out_v[190] = 10'b1011011110;
    16'b0000101100001000: out_v[190] = 10'b1101011010;
    16'b0000100000001000: out_v[190] = 10'b1011100110;
    16'b1000001100000110: out_v[190] = 10'b1000111111;
    16'b0000101000000000: out_v[190] = 10'b0000111110;
    16'b0000000000001000: out_v[190] = 10'b1100011011;
    16'b0000001000100000: out_v[190] = 10'b0110101011;
    16'b0000001000001000: out_v[190] = 10'b0100101101;
    16'b0000101000001000: out_v[190] = 10'b0001110010;
    16'b0000100000101000: out_v[190] = 10'b1000010100;
    16'b0000101000101000: out_v[190] = 10'b0101111011;
    16'b1000100000000000: out_v[190] = 10'b1010100110;
    16'b0000101000100010: out_v[190] = 10'b1000101010;
    16'b0000000000100000: out_v[190] = 10'b0111100100;
    16'b0000101000100000: out_v[190] = 10'b1100010010;
    16'b1000100000000010: out_v[190] = 10'b0111000010;
    16'b0000001000101010: out_v[190] = 10'b1000000100;
    16'b0000000000101000: out_v[190] = 10'b1101011010;
    16'b0000101000101010: out_v[190] = 10'b1000001101;
    16'b0000001000101000: out_v[190] = 10'b1010011011;
    16'b1000100000001000: out_v[190] = 10'b0101101110;
    16'b0000000100001010: out_v[190] = 10'b1101000000;
    16'b0000001100100000: out_v[190] = 10'b1011011111;
    16'b0000000100000010: out_v[190] = 10'b1100110000;
    16'b1000100000001010: out_v[190] = 10'b0010010110;
    16'b0000001100100010: out_v[190] = 10'b0000110010;
    16'b1000101000000010: out_v[190] = 10'b0111001100;
    16'b1000101100000010: out_v[190] = 10'b1011110010;
    16'b0000000000011010: out_v[190] = 10'b0100010110;
    16'b0000000100011000: out_v[190] = 10'b0111001100;
    16'b0000000100011010: out_v[190] = 10'b0111001111;
    16'b0000000000010010: out_v[190] = 10'b1000101001;
    16'b0000000000011000: out_v[190] = 10'b1101100001;
    16'b0000000100010000: out_v[190] = 10'b1001001101;
    16'b0000100000011010: out_v[190] = 10'b0110110011;
    16'b0000000000010000: out_v[190] = 10'b1001001101;
    default: out_v[190] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1000110000000001: out_v[191] = 10'b1001011101;
    16'b1000111000000001: out_v[191] = 10'b1011110111;
    16'b1110111000000001: out_v[191] = 10'b1101011110;
    16'b1110110000000001: out_v[191] = 10'b0010111011;
    16'b0000100000000001: out_v[191] = 10'b1111001010;
    16'b0000111000000001: out_v[191] = 10'b0010100101;
    16'b0110111000000001: out_v[191] = 10'b1100001100;
    16'b0010111000000001: out_v[191] = 10'b0111001100;
    16'b0000011000000001: out_v[191] = 10'b1100100101;
    16'b1000110000000000: out_v[191] = 10'b1001110010;
    16'b1000111000000000: out_v[191] = 10'b1000110111;
    16'b1000110100000001: out_v[191] = 10'b1011001110;
    16'b0000110000000000: out_v[191] = 10'b1101000010;
    16'b1000111100000001: out_v[191] = 10'b0000110011;
    16'b1000110000010001: out_v[191] = 10'b1111011011;
    16'b1000101000000001: out_v[191] = 10'b0101001110;
    16'b0000010000000001: out_v[191] = 10'b1001011101;
    16'b1110100000010001: out_v[191] = 10'b1001101101;
    16'b1000100000000000: out_v[191] = 10'b0101110011;
    16'b1110111000010001: out_v[191] = 10'b1101010011;
    16'b0010110000000001: out_v[191] = 10'b1010010110;
    16'b0110110000000001: out_v[191] = 10'b1110001111;
    16'b1010110000000001: out_v[191] = 10'b0000111110;
    16'b1000111000010001: out_v[191] = 10'b1101001111;
    16'b1000010000000001: out_v[191] = 10'b0000010011;
    16'b1000100000010001: out_v[191] = 10'b1111110110;
    16'b1000011000000001: out_v[191] = 10'b0011100100;
    16'b0000110000000001: out_v[191] = 10'b1000010011;
    16'b1000101000010001: out_v[191] = 10'b1001011110;
    16'b0000100000010001: out_v[191] = 10'b0100011101;
    16'b1010111000000001: out_v[191] = 10'b0111110111;
    16'b1000111100000000: out_v[191] = 10'b1100101101;
    16'b0000011000000000: out_v[191] = 10'b0010101100;
    16'b0000111000000000: out_v[191] = 10'b0110001011;
    16'b1000100000000001: out_v[191] = 10'b0001011111;
    16'b1000101000000000: out_v[191] = 10'b1001001101;
    16'b1000011000000000: out_v[191] = 10'b0111000011;
    16'b0000101000010000: out_v[191] = 10'b1111010011;
    16'b1000010000000000: out_v[191] = 10'b0101100100;
    16'b1010100000000001: out_v[191] = 10'b1111100011;
    16'b1010100000010001: out_v[191] = 10'b1101010111;
    16'b1010110000000000: out_v[191] = 10'b0111111010;
    16'b0110100000010001: out_v[191] = 10'b0100111011;
    16'b0000111000010000: out_v[191] = 10'b1010001001;
    16'b1000001100000000: out_v[191] = 10'b0100011011;
    16'b0000010100000000: out_v[191] = 10'b1001000010;
    16'b0000110100000000: out_v[191] = 10'b1001100010;
    16'b0000010000000000: out_v[191] = 10'b1101101010;
    16'b0000001100000000: out_v[191] = 10'b1001101110;
    16'b0000000100000000: out_v[191] = 10'b0011110101;
    16'b1000001100000001: out_v[191] = 10'b1001101110;
    16'b1000011100000000: out_v[191] = 10'b1110010011;
    16'b0000110100010000: out_v[191] = 10'b1000100110;
    16'b0000011100000000: out_v[191] = 10'b1100110100;
    16'b0000001100000001: out_v[191] = 10'b0110101010;
    16'b1000000100000000: out_v[191] = 10'b1101110011;
    16'b1000010100000000: out_v[191] = 10'b1101100010;
    16'b0000000000000000: out_v[191] = 10'b1101110100;
    16'b0000010100010000: out_v[191] = 10'b1110001001;
    16'b0000101100010000: out_v[191] = 10'b0010111100;
    16'b0000111100010000: out_v[191] = 10'b0100110101;
    16'b0000100100010000: out_v[191] = 10'b0000110101;
    16'b1000101100010000: out_v[191] = 10'b0010011101;
    16'b0000001000000000: out_v[191] = 10'b1010011001;
    16'b0000101000000000: out_v[191] = 10'b1000001011;
    16'b0000001100010000: out_v[191] = 10'b0011001100;
    16'b0000100100000001: out_v[191] = 10'b0100000101;
    16'b0000011100000001: out_v[191] = 10'b1010001000;
    16'b1000001100010000: out_v[191] = 10'b1111001111;
    16'b1000101100000000: out_v[191] = 10'b0111011000;
    16'b0000111100000001: out_v[191] = 10'b1110101000;
    16'b0000010100000001: out_v[191] = 10'b1001011010;
    16'b0000101100010001: out_v[191] = 10'b0011100110;
    16'b1000100100010001: out_v[191] = 10'b0001011111;
    16'b1000101000010000: out_v[191] = 10'b0101111001;
    16'b0000101100000000: out_v[191] = 10'b1101011010;
    16'b0000111100000000: out_v[191] = 10'b1101111001;
    16'b0000000000010001: out_v[191] = 10'b1000011111;
    16'b0000100100010001: out_v[191] = 10'b1100010101;
    16'b0000001000010000: out_v[191] = 10'b0110010101;
    16'b0000101000010001: out_v[191] = 10'b0101110100;
    16'b0000100000000000: out_v[191] = 10'b1001111000;
    16'b1000000000010001: out_v[191] = 10'b1011000110;
    16'b0000000100000001: out_v[191] = 10'b1100001101;
    16'b0000100000010000: out_v[191] = 10'b0011100010;
    16'b0000110100000001: out_v[191] = 10'b0100011111;
    16'b0000000100010001: out_v[191] = 10'b1001011101;
    16'b0000100100000000: out_v[191] = 10'b0111100000;
    16'b1000001000010000: out_v[191] = 10'b0111010000;
    16'b1000000100010001: out_v[191] = 10'b1001011100;
    16'b1000101100010001: out_v[191] = 10'b1011001011;
    16'b0000000100010000: out_v[191] = 10'b0000111101;
    16'b0000000000000001: out_v[191] = 10'b1110001101;
    16'b1000111100010000: out_v[191] = 10'b1001001000;
    16'b1000100000010000: out_v[191] = 10'b0001110100;
    16'b1000101100000001: out_v[191] = 10'b1110010011;
    16'b1000110000010000: out_v[191] = 10'b0111011100;
    16'b1000110100010000: out_v[191] = 10'b1101001101;
    16'b1000100100010000: out_v[191] = 10'b0011110011;
    16'b1000111000010000: out_v[191] = 10'b1101011111;
    16'b1000000100000001: out_v[191] = 10'b1110101110;
    16'b1000111100010001: out_v[191] = 10'b0010100010;
    16'b1000100100000001: out_v[191] = 10'b1110010010;
    16'b0000110000010000: out_v[191] = 10'b1010001001;
    16'b1000110100000000: out_v[191] = 10'b0110110010;
    16'b1000100100000000: out_v[191] = 10'b0110110100;
    16'b1000010100000001: out_v[191] = 10'b0101010011;
    16'b0110100100000001: out_v[191] = 10'b0010100110;
    16'b0110101100000000: out_v[191] = 10'b0000110011;
    16'b1000011100000001: out_v[191] = 10'b1110101101;
    16'b0000101100000001: out_v[191] = 10'b0100110010;
    16'b0010100100000001: out_v[191] = 10'b0001110110;
    16'b0010101100000000: out_v[191] = 10'b0100110011;
    16'b0110100000000001: out_v[191] = 10'b1011101111;
    16'b1000000000000001: out_v[191] = 10'b1010001010;
    16'b0010000100000001: out_v[191] = 10'b0101011111;
    16'b1000000100010000: out_v[191] = 10'b1000111001;
    16'b1000000000000000: out_v[191] = 10'b0101110101;
    16'b1000000000010000: out_v[191] = 10'b1011110011;
    16'b0000000000010000: out_v[191] = 10'b0011110100;
    16'b0010100100010000: out_v[191] = 10'b1001001110;
    16'b0000100001010000: out_v[191] = 10'b0111000011;
    16'b0000110101000000: out_v[191] = 10'b0111100101;
    16'b0010100000010000: out_v[191] = 10'b1011001010;
    16'b0000100101010000: out_v[191] = 10'b1101000001;
    16'b1000001000000000: out_v[191] = 10'b0101011011;
    16'b1100011000000001: out_v[191] = 10'b1011100110;
    16'b0000111000001100: out_v[191] = 10'b1011110011;
    16'b0110111000000000: out_v[191] = 10'b1101010111;
    16'b0100111000001100: out_v[191] = 10'b0101110111;
    16'b0000111000001101: out_v[191] = 10'b1111110100;
    16'b0100111000001101: out_v[191] = 10'b1111110111;
    16'b0000011000001101: out_v[191] = 10'b1111001011;
    16'b0000111000001000: out_v[191] = 10'b1011110001;
    16'b0000011000001000: out_v[191] = 10'b1111001001;
    16'b1000011000001101: out_v[191] = 10'b0111100000;
    16'b1110011000000001: out_v[191] = 10'b1000011011;
    16'b0000011000001100: out_v[191] = 10'b1101111001;
    16'b0110111000001101: out_v[191] = 10'b0110001111;
    16'b1000011000001001: out_v[191] = 10'b1101111001;
    16'b1010011000000001: out_v[191] = 10'b0111101011;
    16'b1000110100010001: out_v[191] = 10'b1110100011;
    16'b0110111100000000: out_v[191] = 10'b1001001100;
    16'b0010111100000000: out_v[191] = 10'b0100010001;
    16'b0110111100000001: out_v[191] = 10'b1100000101;
    16'b0010111100000001: out_v[191] = 10'b1001101011;
    default: out_v[191] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000001110010: out_v[192] = 10'b0100011111;
    16'b0100000001010001: out_v[192] = 10'b1001100001;
    16'b0100000000000011: out_v[192] = 10'b1100000101;
    16'b0100000000110011: out_v[192] = 10'b0110000001;
    16'b0100000001110000: out_v[192] = 10'b0011010011;
    16'b0000000001100011: out_v[192] = 10'b0010101101;
    16'b0000000001110011: out_v[192] = 10'b0110001101;
    16'b0100000000000010: out_v[192] = 10'b0011111101;
    16'b0000000000110010: out_v[192] = 10'b0111011010;
    16'b0100000001110001: out_v[192] = 10'b1111100001;
    16'b0000000001110000: out_v[192] = 10'b1000001011;
    16'b0100000000010011: out_v[192] = 10'b1111000010;
    16'b0000000000000011: out_v[192] = 10'b0111111001;
    16'b0000000001010001: out_v[192] = 10'b0010110100;
    16'b0100000000100011: out_v[192] = 10'b0000000101;
    16'b0100000001110011: out_v[192] = 10'b0100001001;
    16'b0000000000010011: out_v[192] = 10'b1000011110;
    16'b0100000000110010: out_v[192] = 10'b0101011010;
    16'b0000000000100011: out_v[192] = 10'b0101010100;
    16'b0100000000100010: out_v[192] = 10'b0000000111;
    16'b0000000001000011: out_v[192] = 10'b0011001011;
    16'b0100000001000011: out_v[192] = 10'b1111011011;
    16'b0000000000110011: out_v[192] = 10'b0111011011;
    16'b0100000001010011: out_v[192] = 10'b1011000001;
    16'b0000000001010000: out_v[192] = 10'b0000110110;
    16'b0100000001010000: out_v[192] = 10'b0101110001;
    16'b0000000000100010: out_v[192] = 10'b1110110100;
    16'b0000000000000010: out_v[192] = 10'b0010101011;
    16'b0100000001010010: out_v[192] = 10'b1000010110;
    16'b0000000001010011: out_v[192] = 10'b1010101010;
    16'b0100000000010010: out_v[192] = 10'b0000100101;
    16'b0000000000010010: out_v[192] = 10'b0001110110;
    16'b0000000000100001: out_v[192] = 10'b0111100011;
    16'b0000000001110001: out_v[192] = 10'b1101011010;
    16'b0100000001110010: out_v[192] = 10'b1110111100;
    16'b0000000001100010: out_v[192] = 10'b1110011101;
    16'b0100000001100000: out_v[192] = 10'b0100011011;
    16'b0000000001000000: out_v[192] = 10'b0011001010;
    16'b0000000001000010: out_v[192] = 10'b0100111010;
    16'b0100000000100000: out_v[192] = 10'b1100011111;
    16'b0000000001100000: out_v[192] = 10'b0010101110;
    16'b0100000001000000: out_v[192] = 10'b1000101010;
    16'b0000000000100000: out_v[192] = 10'b1101010101;
    16'b0000000000000000: out_v[192] = 10'b1101001100;
    16'b0100000000000000: out_v[192] = 10'b0100100011;
    16'b0000000000110000: out_v[192] = 10'b1101110101;
    16'b0100000001100011: out_v[192] = 10'b1001010110;
    16'b0100000000000001: out_v[192] = 10'b0001101111;
    16'b0100000001100010: out_v[192] = 10'b1100110100;
    16'b0000000000010000: out_v[192] = 10'b1100011100;
    16'b0000000001100001: out_v[192] = 10'b0101001110;
    16'b0100000000100001: out_v[192] = 10'b0000011110;
    16'b0100000000110000: out_v[192] = 10'b1100101010;
    16'b0100000001100001: out_v[192] = 10'b0110110100;
    16'b0000000001010010: out_v[192] = 10'b1110001110;
    16'b0100000000010000: out_v[192] = 10'b1000101000;
    16'b0100000001000010: out_v[192] = 10'b0001001010;
    16'b0000000000000001: out_v[192] = 10'b1010000001;
    16'b0000000000010001: out_v[192] = 10'b1010000010;
    16'b0000000000110001: out_v[192] = 10'b1111100011;
    16'b0010000000100001: out_v[192] = 10'b0111100011;
    16'b0010000000110000: out_v[192] = 10'b1111101011;
    16'b0000000001000001: out_v[192] = 10'b1011000010;
    16'b0000000011000000: out_v[192] = 10'b1101111110;
    default: out_v[192] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010001000000000: out_v[193] = 10'b0000011111;
    16'b0000001000000000: out_v[193] = 10'b0010010100;
    16'b0010101000000000: out_v[193] = 10'b1000001011;
    16'b0111001000000000: out_v[193] = 10'b1001001000;
    16'b0011001000000000: out_v[193] = 10'b1001100100;
    16'b0001001000000000: out_v[193] = 10'b0101000101;
    16'b0010100000000010: out_v[193] = 10'b1111110101;
    16'b0000100000000000: out_v[193] = 10'b1110001001;
    16'b0000000000000000: out_v[193] = 10'b1010001011;
    16'b0010001000000010: out_v[193] = 10'b1000010101;
    16'b0000101000000000: out_v[193] = 10'b0111000011;
    16'b0011101000010100: out_v[193] = 10'b1100100101;
    16'b0000100000010100: out_v[193] = 10'b0010011010;
    16'b0100000000000000: out_v[193] = 10'b0001010111;
    16'b0010000000000000: out_v[193] = 10'b1110111011;
    16'b0100101000000000: out_v[193] = 10'b0001110011;
    16'b0010101000000010: out_v[193] = 10'b1010110111;
    16'b0011001000000010: out_v[193] = 10'b1101110010;
    16'b0011101000000000: out_v[193] = 10'b0011101011;
    16'b0010101000000011: out_v[193] = 10'b1001011010;
    16'b0000001000000011: out_v[193] = 10'b1011011011;
    16'b0010000000000010: out_v[193] = 10'b0001101111;
    16'b0010001000000011: out_v[193] = 10'b0011000111;
    16'b0100100000000000: out_v[193] = 10'b0001111110;
    16'b0100001000000000: out_v[193] = 10'b0101010000;
    16'b0001101000010100: out_v[193] = 10'b1001011111;
    16'b0110001000000000: out_v[193] = 10'b0000111010;
    16'b0110101000000000: out_v[193] = 10'b1100101110;
    16'b0010100000000000: out_v[193] = 10'b1011100111;
    16'b0001001000010100: out_v[193] = 10'b0011101000;
    16'b0001101000000000: out_v[193] = 10'b1101101100;
    16'b0000001000010100: out_v[193] = 10'b1000110110;
    16'b0001001000000100: out_v[193] = 10'b1110100001;
    16'b0010000000000011: out_v[193] = 10'b1000010101;
    16'b0010001000010100: out_v[193] = 10'b1010100000;
    16'b0000101000010100: out_v[193] = 10'b1000111101;
    16'b0010101000010100: out_v[193] = 10'b1101001011;
    16'b0011001000010100: out_v[193] = 10'b1110111001;
    16'b0101001000000000: out_v[193] = 10'b1100100010;
    16'b0111101000000000: out_v[193] = 10'b1111000011;
    16'b0000101000000100: out_v[193] = 10'b0011101110;
    16'b0000000000010100: out_v[193] = 10'b0100011001;
    16'b0001100000010100: out_v[193] = 10'b1100010011;
    16'b0001100000000000: out_v[193] = 10'b0000111010;
    16'b0000100000000100: out_v[193] = 10'b1111100001;
    16'b0001101000000100: out_v[193] = 10'b1010110111;
    16'b0000000000000100: out_v[193] = 10'b1100100110;
    16'b0001100000000100: out_v[193] = 10'b1001110011;
    16'b0010101000010111: out_v[193] = 10'b1111011000;
    16'b0010101000000001: out_v[193] = 10'b1001010100;
    16'b0001000000000000: out_v[193] = 10'b1011000101;
    16'b0010100000000001: out_v[193] = 10'b1011100100;
    16'b0011100000010111: out_v[193] = 10'b1000111110;
    16'b0010100000010111: out_v[193] = 10'b1111010111;
    16'b0010100000010100: out_v[193] = 10'b0101110100;
    16'b0011000000000000: out_v[193] = 10'b1110100001;
    16'b0111000000000001: out_v[193] = 10'b1001001111;
    16'b0111000000010100: out_v[193] = 10'b1011110111;
    16'b0010000000000001: out_v[193] = 10'b1101100110;
    16'b0000000000010110: out_v[193] = 10'b1111011100;
    16'b0000100000000010: out_v[193] = 10'b1001010101;
    16'b0010100000000011: out_v[193] = 10'b0001111011;
    16'b0011000000000001: out_v[193] = 10'b1111111011;
    16'b0010000000010100: out_v[193] = 10'b0110101010;
    16'b0010101000010110: out_v[193] = 10'b1000001101;
    16'b0111000000000000: out_v[193] = 10'b1111100110;
    16'b0010100000010110: out_v[193] = 10'b1101011110;
    16'b0011000000010100: out_v[193] = 10'b0101001101;
    16'b0000100000010110: out_v[193] = 10'b0011000100;
    16'b0000000000000010: out_v[193] = 10'b1101001111;
    16'b0011101000010111: out_v[193] = 10'b1100010111;
    16'b0010100000010101: out_v[193] = 10'b0011010101;
    16'b0011001000000001: out_v[193] = 10'b0011011100;
    16'b0101000000000000: out_v[193] = 10'b1011100001;
    16'b0001000000010100: out_v[193] = 10'b0111010100;
    16'b0010001000000001: out_v[193] = 10'b1111110110;
    16'b0011101000010110: out_v[193] = 10'b1110011111;
    16'b0101101000000000: out_v[193] = 10'b0101110010;
    16'b0010101000000100: out_v[193] = 10'b0101011110;
    16'b0110101000010100: out_v[193] = 10'b0010111111;
    16'b0101101000010100: out_v[193] = 10'b0111010010;
    16'b0100001000010100: out_v[193] = 10'b0101011011;
    16'b0010100000000100: out_v[193] = 10'b0101101011;
    16'b0111101000010100: out_v[193] = 10'b1111101001;
    16'b0010000000000100: out_v[193] = 10'b1111101111;
    16'b0000001000000100: out_v[193] = 10'b0110010011;
    16'b0000101001010100: out_v[193] = 10'b1000111110;
    16'b0010001001010100: out_v[193] = 10'b1001001100;
    16'b0010001000010111: out_v[193] = 10'b0000110110;
    16'b0010001000000100: out_v[193] = 10'b1010100011;
    16'b0000001001010100: out_v[193] = 10'b1011011111;
    16'b0011000100000000: out_v[193] = 10'b0001011001;
    16'b0010000000010110: out_v[193] = 10'b1000011000;
    16'b0000000100010100: out_v[193] = 10'b1111001011;
    16'b0001000000000100: out_v[193] = 10'b1110011101;
    16'b0010000100000000: out_v[193] = 10'b1110101010;
    16'b0000000100000000: out_v[193] = 10'b0001010010;
    16'b0011000100010100: out_v[193] = 10'b0110010101;
    16'b0010000100000010: out_v[193] = 10'b0011111111;
    16'b0001000100000000: out_v[193] = 10'b0111101011;
    16'b0001000100010100: out_v[193] = 10'b0011011111;
    16'b0010000100010100: out_v[193] = 10'b1111101010;
    16'b0010000100000100: out_v[193] = 10'b1011111101;
    16'b0001000000100000: out_v[193] = 10'b1011101011;
    16'b0000000100000100: out_v[193] = 10'b0101111011;
    16'b0011000000000100: out_v[193] = 10'b1001011111;
    16'b0000101000001000: out_v[193] = 10'b0111000001;
    16'b0000001000001000: out_v[193] = 10'b0010111011;
    16'b0000100000001000: out_v[193] = 10'b1010100100;
    16'b0000000000001000: out_v[193] = 10'b0011010101;
    16'b0000001000011100: out_v[193] = 10'b1001000111;
    16'b0000101000011100: out_v[193] = 10'b1001010111;
    default: out_v[193] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1011000000100000: out_v[194] = 10'b1101000100;
    16'b1001000000000001: out_v[194] = 10'b0110101000;
    16'b1011010000010101: out_v[194] = 10'b1110110011;
    16'b1011000000000000: out_v[194] = 10'b1010011001;
    16'b0011011000010101: out_v[194] = 10'b0000011111;
    16'b1011000000000001: out_v[194] = 10'b0011100011;
    16'b0001011000010101: out_v[194] = 10'b1011100011;
    16'b1001000000100000: out_v[194] = 10'b1001010001;
    16'b0011000000010101: out_v[194] = 10'b0111011011;
    16'b0001000000000001: out_v[194] = 10'b1101111100;
    16'b0011000000000101: out_v[194] = 10'b1011111100;
    16'b1001000000000000: out_v[194] = 10'b0011101100;
    16'b0011000000000000: out_v[194] = 10'b0000101000;
    16'b0010000000010101: out_v[194] = 10'b0010001011;
    16'b0011010000010101: out_v[194] = 10'b1110111110;
    16'b0010010000010101: out_v[194] = 10'b0011011111;
    16'b0010011000010101: out_v[194] = 10'b0110001110;
    16'b1011011000110101: out_v[194] = 10'b0010001011;
    16'b0000011000010101: out_v[194] = 10'b0100100001;
    16'b1011000000000101: out_v[194] = 10'b0011010101;
    16'b0011011000110101: out_v[194] = 10'b0011000011;
    16'b1001000000100001: out_v[194] = 10'b1000111100;
    16'b0001010000010101: out_v[194] = 10'b0001111111;
    16'b0010000000000100: out_v[194] = 10'b1100001011;
    16'b0011000000000001: out_v[194] = 10'b0111000111;
    16'b1000000000000001: out_v[194] = 10'b0000110111;
    16'b1011010000000001: out_v[194] = 10'b1110000111;
    16'b0001000000000000: out_v[194] = 10'b0110111010;
    16'b0001000000000101: out_v[194] = 10'b0100111111;
    16'b0011000000000100: out_v[194] = 10'b1011110100;
    16'b0001011000000001: out_v[194] = 10'b0011010011;
    16'b0010000000010100: out_v[194] = 10'b0110001111;
    16'b1011010000110101: out_v[194] = 10'b0011111011;
    16'b0000010000010101: out_v[194] = 10'b0010111110;
    16'b1011010000000101: out_v[194] = 10'b0100111111;
    16'b1011000000100001: out_v[194] = 10'b1000101010;
    16'b0011010000110101: out_v[194] = 10'b0011100111;
    16'b0000000000100000: out_v[194] = 10'b0000101110;
    16'b0000000000000000: out_v[194] = 10'b1010001101;
    16'b0010000000100000: out_v[194] = 10'b0010111010;
    16'b0000000000100010: out_v[194] = 10'b1110101010;
    16'b0001000000100000: out_v[194] = 10'b1101000100;
    16'b0001000000100100: out_v[194] = 10'b1011110100;
    16'b1001000000010101: out_v[194] = 10'b1111100110;
    16'b0001000000110100: out_v[194] = 10'b1000011100;
    16'b0000000000100100: out_v[194] = 10'b1011011011;
    16'b0001000000000100: out_v[194] = 10'b1010110010;
    16'b1001000000100100: out_v[194] = 10'b0111100111;
    16'b0000000000110100: out_v[194] = 10'b1111100110;
    16'b1000000000010101: out_v[194] = 10'b0001101011;
    16'b0011000000110100: out_v[194] = 10'b1000100110;
    16'b1001000000000100: out_v[194] = 10'b0011101111;
    16'b1010000000100001: out_v[194] = 10'b1000100111;
    16'b1000000000100000: out_v[194] = 10'b0101000000;
    16'b1010000000100101: out_v[194] = 10'b1011100110;
    16'b0001000000010100: out_v[194] = 10'b0110010010;
    16'b1000000000010100: out_v[194] = 10'b0000101011;
    16'b1011000000110101: out_v[194] = 10'b1100110110;
    16'b0001000000100101: out_v[194] = 10'b0000110101;
    16'b1011000000110100: out_v[194] = 10'b0000010101;
    16'b0001010000110100: out_v[194] = 10'b0010110111;
    16'b1000010000110100: out_v[194] = 10'b0101010111;
    16'b1010000000100000: out_v[194] = 10'b0110011010;
    16'b1001000000110100: out_v[194] = 10'b0111000010;
    16'b0001000000110101: out_v[194] = 10'b1010110011;
    16'b1000000000100001: out_v[194] = 10'b1101100011;
    16'b1000000000100100: out_v[194] = 10'b1100110110;
    16'b0001000000100001: out_v[194] = 10'b1000100101;
    16'b0011000000100001: out_v[194] = 10'b1000111101;
    16'b1010000000110101: out_v[194] = 10'b1110111000;
    16'b1000000000000100: out_v[194] = 10'b0001111010;
    16'b1011000000100100: out_v[194] = 10'b0101100110;
    16'b0011000000100000: out_v[194] = 10'b0101101100;
    16'b1000000000110101: out_v[194] = 10'b1000011111;
    16'b1010000000000101: out_v[194] = 10'b0111110111;
    16'b1001010000110100: out_v[194] = 10'b1111100000;
    16'b1011000000100101: out_v[194] = 10'b1011011000;
    16'b1000000000110100: out_v[194] = 10'b1101001011;
    16'b0011000000100100: out_v[194] = 10'b1000000101;
    16'b1000010000100000: out_v[194] = 10'b0100100111;
    16'b1011000000010101: out_v[194] = 10'b0011000110;
    16'b1000010000110000: out_v[194] = 10'b1101001001;
    16'b1001000000010100: out_v[194] = 10'b1001001101;
    16'b1000000000000000: out_v[194] = 10'b0010111000;
    16'b1010000000000000: out_v[194] = 10'b1010001011;
    16'b0001010000010100: out_v[194] = 10'b1000111100;
    16'b0000010000010100: out_v[194] = 10'b1111111000;
    16'b0000000000000100: out_v[194] = 10'b1100110000;
    16'b0000000000010100: out_v[194] = 10'b1000011110;
    16'b1011000000000100: out_v[194] = 10'b0011001110;
    16'b1001010000010100: out_v[194] = 10'b1011100001;
    16'b0000000000000001: out_v[194] = 10'b0010100011;
    16'b1000010000000001: out_v[194] = 10'b0101011110;
    16'b0010000000000000: out_v[194] = 10'b1010000101;
    16'b1010000000000001: out_v[194] = 10'b1010001010;
    16'b1000000000000101: out_v[194] = 10'b0000111100;
    16'b1001010000000001: out_v[194] = 10'b0111101011;
    16'b0010000000000001: out_v[194] = 10'b0010011011;
    16'b1001000000000010: out_v[194] = 10'b0001110010;
    16'b0001000000000010: out_v[194] = 10'b0001010010;
    16'b1101000000100000: out_v[194] = 10'b0100011111;
    16'b1001011000110101: out_v[194] = 10'b0011111011;
    16'b0001011000110100: out_v[194] = 10'b1111011010;
    16'b1001010000110101: out_v[194] = 10'b1101001010;
    16'b0001011000110101: out_v[194] = 10'b0011011111;
    16'b1101000000000000: out_v[194] = 10'b1101110100;
    16'b1101000000100001: out_v[194] = 10'b1111100011;
    16'b0101000000100000: out_v[194] = 10'b1111100101;
    16'b0001010000110101: out_v[194] = 10'b0101000111;
    16'b1010000000100100: out_v[194] = 10'b1101011011;
    default: out_v[194] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000000000010: out_v[195] = 10'b1011100101;
    16'b0000000010000110: out_v[195] = 10'b0001000001;
    16'b0001000010000110: out_v[195] = 10'b1101010101;
    16'b0000000000000100: out_v[195] = 10'b1110010001;
    16'b0000000000000110: out_v[195] = 10'b0111001011;
    16'b0001000010000100: out_v[195] = 10'b0100010101;
    16'b0000000000000000: out_v[195] = 10'b1110110110;
    16'b0000000001000110: out_v[195] = 10'b0101101010;
    16'b0000000010000100: out_v[195] = 10'b0100010011;
    16'b0000000010000010: out_v[195] = 10'b0011000100;
    16'b0000000010000000: out_v[195] = 10'b0110110101;
    16'b0000000011000110: out_v[195] = 10'b0101111010;
    16'b0001000011000100: out_v[195] = 10'b0010100111;
    16'b0000000011000100: out_v[195] = 10'b1011110100;
    16'b0000000001000000: out_v[195] = 10'b1110000111;
    16'b0000000001000010: out_v[195] = 10'b0110001010;
    16'b0000000011000000: out_v[195] = 10'b1100010011;
    16'b0000000001000100: out_v[195] = 10'b1001000110;
    16'b0000000011000010: out_v[195] = 10'b1100101010;
    16'b0001000010000000: out_v[195] = 10'b0001001100;
    16'b0001000001000100: out_v[195] = 10'b1111000110;
    16'b0000000001000001: out_v[195] = 10'b0100011100;
    16'b0000000001000011: out_v[195] = 10'b0110000010;
    16'b0001000001000000: out_v[195] = 10'b1000101010;
    16'b0000000000000001: out_v[195] = 10'b0010001011;
    16'b0001000011000000: out_v[195] = 10'b0110001010;
    16'b0000000000000011: out_v[195] = 10'b1011000110;
    16'b0001000000000000: out_v[195] = 10'b0110110111;
    16'b0001000000000100: out_v[195] = 10'b1111010000;
    16'b0001000001000010: out_v[195] = 10'b0001001001;
    16'b0001000011000010: out_v[195] = 10'b0011111000;
    16'b0000000001000111: out_v[195] = 10'b1011101000;
    16'b0000000000000101: out_v[195] = 10'b0110010111;
    16'b0000000001000101: out_v[195] = 10'b0011101000;
    16'b0000000010001000: out_v[195] = 10'b0010111010;
    16'b0000000011001010: out_v[195] = 10'b1000100110;
    16'b0000000010001010: out_v[195] = 10'b1101111001;
    16'b0000000011001000: out_v[195] = 10'b1011001100;
    16'b1000000000000100: out_v[195] = 10'b1011001100;
    16'b1000000001000000: out_v[195] = 10'b1100111001;
    16'b1000000000000000: out_v[195] = 10'b1101000110;
    16'b1000000001000100: out_v[195] = 10'b0101000101;
    16'b0000001000000010: out_v[195] = 10'b0010010010;
    16'b0000001000000000: out_v[195] = 10'b0001010001;
    default: out_v[195] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000010000010: out_v[196] = 10'b1101000011;
    16'b0000010010000000: out_v[196] = 10'b0110011110;
    16'b0000000010000110: out_v[196] = 10'b1100001011;
    16'b0000010010000110: out_v[196] = 10'b1111001100;
    16'b0000000010000000: out_v[196] = 10'b1110000011;
    16'b0000100010000000: out_v[196] = 10'b1000010011;
    16'b0000000010000100: out_v[196] = 10'b1000011011;
    16'b0000000000000100: out_v[196] = 10'b1111000111;
    16'b0000000000000000: out_v[196] = 10'b1111100010;
    16'b0000000000000010: out_v[196] = 10'b0011100010;
    16'b0000100010000110: out_v[196] = 10'b1110010011;
    16'b0000010000000100: out_v[196] = 10'b0001001011;
    16'b0000010000000000: out_v[196] = 10'b0001101011;
    16'b0000000000000110: out_v[196] = 10'b0010111000;
    16'b0000110010000100: out_v[196] = 10'b0110001111;
    16'b0000010000000110: out_v[196] = 10'b1000010111;
    16'b0000110000000100: out_v[196] = 10'b1101110111;
    16'b0000010010000100: out_v[196] = 10'b0100011000;
    16'b0000100010000010: out_v[196] = 10'b0011110010;
    16'b0000110010000000: out_v[196] = 10'b0110010111;
    16'b0100100110000000: out_v[196] = 10'b0111000010;
    16'b0100100100000000: out_v[196] = 10'b1011111101;
    16'b0100000100000000: out_v[196] = 10'b1001110010;
    16'b0100000000000000: out_v[196] = 10'b1110100100;
    16'b0100000010000000: out_v[196] = 10'b0111011010;
    16'b0100000110000000: out_v[196] = 10'b1010110110;
    16'b0100110110000000: out_v[196] = 10'b1111100011;
    16'b0100000000000010: out_v[196] = 10'b0010101010;
    16'b0100100110000010: out_v[196] = 10'b1001001000;
    16'b0100100111000010: out_v[196] = 10'b1111000100;
    16'b0100100011000000: out_v[196] = 10'b0110011111;
    16'b0000100110000010: out_v[196] = 10'b0010011011;
    16'b0100100000000000: out_v[196] = 10'b1100011011;
    16'b0100100100000010: out_v[196] = 10'b1111011001;
    16'b0000100110000000: out_v[196] = 10'b1010111000;
    16'b0100110110000100: out_v[196] = 10'b1010101101;
    16'b0100100010000100: out_v[196] = 10'b0111100110;
    16'b0100000010000010: out_v[196] = 10'b0011001010;
    16'b0100100010000000: out_v[196] = 10'b0100001101;
    16'b0100110110000010: out_v[196] = 10'b0010111100;
    16'b0000110110000010: out_v[196] = 10'b1000100011;
    16'b0100100110000110: out_v[196] = 10'b1001001000;
    16'b0000100100000000: out_v[196] = 10'b0001111100;
    16'b0100110010000000: out_v[196] = 10'b1111001011;
    16'b0100100111000000: out_v[196] = 10'b1010100111;
    16'b0000100100000010: out_v[196] = 10'b0111000111;
    16'b0100110110000110: out_v[196] = 10'b1010010010;
    16'b0100000010000100: out_v[196] = 10'b0010110100;
    16'b0100100010000110: out_v[196] = 10'b0011011111;
    16'b0100100110000100: out_v[196] = 10'b1011001100;
    16'b0000100000000010: out_v[196] = 10'b0011100101;
    16'b0100100010000010: out_v[196] = 10'b0110010111;
    16'b0000100111000010: out_v[196] = 10'b0101101001;
    16'b0100000011000010: out_v[196] = 10'b1010110011;
    16'b0100000011000000: out_v[196] = 10'b1011111010;
    16'b0000110110000000: out_v[196] = 10'b1010100110;
    16'b0100110010000100: out_v[196] = 10'b1011101101;
    16'b0100010000000100: out_v[196] = 10'b0011010111;
    16'b0100110000000000: out_v[196] = 10'b1101101000;
    16'b0100010010000000: out_v[196] = 10'b0000010101;
    16'b0000110010000010: out_v[196] = 10'b1111010101;
    16'b0000100000000000: out_v[196] = 10'b0110001100;
    16'b0000110100000010: out_v[196] = 10'b0000010010;
    16'b0000110100000000: out_v[196] = 10'b1000110000;
    16'b0000110000000000: out_v[196] = 10'b0011100100;
    16'b0100100000000010: out_v[196] = 10'b0100011010;
    16'b0100110100000010: out_v[196] = 10'b1010001011;
    16'b0100110100000000: out_v[196] = 10'b0100001010;
    16'b0000100110000110: out_v[196] = 10'b1110111011;
    16'b0100010000000000: out_v[196] = 10'b1010110111;
    16'b0000110000000010: out_v[196] = 10'b1100110110;
    16'b0000100110000100: out_v[196] = 10'b0001111010;
    16'b0100010000000010: out_v[196] = 10'b1011010010;
    16'b0100100100000100: out_v[196] = 10'b1110011100;
    16'b0100100000000100: out_v[196] = 10'b1100010110;
    16'b0100100000000110: out_v[196] = 10'b0001111001;
    16'b0100100100000110: out_v[196] = 10'b0100011100;
    16'b0100000000000100: out_v[196] = 10'b0000110110;
    16'b0100100101000010: out_v[196] = 10'b1111000010;
    16'b0000100111000000: out_v[196] = 10'b0001011100;
    16'b0000100011000000: out_v[196] = 10'b0011011110;
    16'b0100100101000000: out_v[196] = 10'b0001000001;
    16'b0000101000000000: out_v[196] = 10'b0110010011;
    16'b0100000100000010: out_v[196] = 10'b1101000101;
    default: out_v[196] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000000000000: out_v[197] = 10'b1000100010;
    16'b0000000000010010: out_v[197] = 10'b1011000101;
    16'b0000000001010010: out_v[197] = 10'b1101100110;
    16'b0000001001010010: out_v[197] = 10'b1100111111;
    16'b0000000001000010: out_v[197] = 10'b0010011101;
    16'b0000000000011010: out_v[197] = 10'b0101011100;
    16'b0000000011010010: out_v[197] = 10'b1111000011;
    16'b0000000000000010: out_v[197] = 10'b1110110011;
    16'b0000000000001010: out_v[197] = 10'b1111111001;
    16'b0110001011010000: out_v[197] = 10'b1000101011;
    16'b0000000000010000: out_v[197] = 10'b0011001011;
    16'b0000000000011110: out_v[197] = 10'b0010110010;
    16'b0000000000011100: out_v[197] = 10'b1101100100;
    16'b0100000001010010: out_v[197] = 10'b0011110011;
    16'b0000001000010010: out_v[197] = 10'b0111010011;
    16'b0000000010010010: out_v[197] = 10'b0111100000;
    16'b0100001001010010: out_v[197] = 10'b0111110101;
    16'b0110000011011010: out_v[197] = 10'b1001001010;
    16'b0000000000011000: out_v[197] = 10'b1001000110;
    16'b0100000011010010: out_v[197] = 10'b0100111111;
    16'b0100001011010010: out_v[197] = 10'b1010111101;
    16'b0100001001011010: out_v[197] = 10'b1110001011;
    16'b0010000011010000: out_v[197] = 10'b1011011111;
    16'b0000001000011010: out_v[197] = 10'b0110010101;
    16'b0110000011010010: out_v[197] = 10'b1111001011;
    16'b0110001011010010: out_v[197] = 10'b1011010110;
    16'b0000000000001000: out_v[197] = 10'b1110110110;
    16'b0000000001011010: out_v[197] = 10'b1010101111;
    16'b0000000000010110: out_v[197] = 10'b0011001100;
    16'b0000000010011010: out_v[197] = 10'b0111001110;
    16'b0110000011010000: out_v[197] = 10'b1101011100;
    16'b0000001001011010: out_v[197] = 10'b1110110111;
    16'b0100000011011010: out_v[197] = 10'b1011011010;
    16'b0000000000010100: out_v[197] = 10'b0101010111;
    16'b0110001011011010: out_v[197] = 10'b1111010110;
    16'b0100001011011010: out_v[197] = 10'b0110101110;
    16'b0000000010000010: out_v[197] = 10'b0011111110;
    16'b0100000001011010: out_v[197] = 10'b1111100010;
    16'b0000000011011010: out_v[197] = 10'b1001110110;
    16'b0000000000001100: out_v[197] = 10'b1101011111;
    16'b0000001000001000: out_v[197] = 10'b1101011000;
    16'b0000000000000100: out_v[197] = 10'b1000010010;
    16'b0000001000000000: out_v[197] = 10'b1010001111;
    16'b0000001000001100: out_v[197] = 10'b0001100011;
    16'b0000001000000100: out_v[197] = 10'b1101011100;
    16'b0100001000001100: out_v[197] = 10'b1111000110;
    16'b0110001011001100: out_v[197] = 10'b1011011101;
    16'b0000001000011110: out_v[197] = 10'b1010110110;
    16'b0000001010011100: out_v[197] = 10'b1110111110;
    16'b0110000011001101: out_v[197] = 10'b1110100100;
    16'b0000000001001100: out_v[197] = 10'b0110010100;
    16'b0010001010011100: out_v[197] = 10'b1101111101;
    16'b0000001000011000: out_v[197] = 10'b1010111011;
    16'b0000001000011100: out_v[197] = 10'b0011101110;
    16'b0100001011011100: out_v[197] = 10'b1011100001;
    16'b0110001011011000: out_v[197] = 10'b0101111111;
    16'b0010000010011100: out_v[197] = 10'b0000011111;
    16'b0010001010011000: out_v[197] = 10'b1110001111;
    16'b0110001011011101: out_v[197] = 10'b0111111001;
    16'b0110001011011100: out_v[197] = 10'b0011111001;
    16'b0100001001001100: out_v[197] = 10'b1000101001;
    16'b0000000010011000: out_v[197] = 10'b1101110100;
    16'b0100001011001100: out_v[197] = 10'b0111011000;
    16'b0100000001011110: out_v[197] = 10'b0000110101;
    16'b0110000011001100: out_v[197] = 10'b1101010101;
    16'b0010001010011110: out_v[197] = 10'b1000110111;
    16'b0110000011011100: out_v[197] = 10'b0000001101;
    16'b0100001011011110: out_v[197] = 10'b1111111010;
    16'b0110001010011100: out_v[197] = 10'b1000010011;
    16'b0110001011011110: out_v[197] = 10'b0111111011;
    16'b0110001011001101: out_v[197] = 10'b1111100111;
    16'b0100001001011100: out_v[197] = 10'b1011101100;
    16'b0100001001011110: out_v[197] = 10'b1011110110;
    16'b0100001001011000: out_v[197] = 10'b0010011110;
    16'b0100000001001100: out_v[197] = 10'b0011110010;
    16'b0100000001000110: out_v[197] = 10'b0000110110;
    16'b0100000001000101: out_v[197] = 10'b1110110111;
    16'b0100000001010100: out_v[197] = 10'b0110111010;
    16'b0100000001000000: out_v[197] = 10'b0000111010;
    16'b0100000001000100: out_v[197] = 10'b1001100011;
    16'b0000000000000110: out_v[197] = 10'b0010101110;
    16'b0000001000000110: out_v[197] = 10'b1001101000;
    16'b0110000011000111: out_v[197] = 10'b1010001000;
    16'b0110000011000011: out_v[197] = 10'b1001101001;
    16'b0100000001000010: out_v[197] = 10'b1011100111;
    16'b0100000001000111: out_v[197] = 10'b0011000011;
    16'b0100001001000110: out_v[197] = 10'b1011001110;
    16'b0000000001000000: out_v[197] = 10'b0011101110;
    16'b0100000011000111: out_v[197] = 10'b1001110011;
    16'b0110000011000110: out_v[197] = 10'b1000111010;
    16'b0000000001000100: out_v[197] = 10'b1010011101;
    16'b0100001001000100: out_v[197] = 10'b0001111011;
    16'b0000001000001110: out_v[197] = 10'b1101011001;
    16'b0100001000000110: out_v[197] = 10'b1101010111;
    16'b0000000001000110: out_v[197] = 10'b0000001110;
    16'b0100000000000100: out_v[197] = 10'b0000001011;
    16'b0000001000010100: out_v[197] = 10'b0110010010;
    16'b0100001000000100: out_v[197] = 10'b1100001010;
    16'b0100000001001110: out_v[197] = 10'b1101010001;
    16'b0100000011000110: out_v[197] = 10'b0010110110;
    16'b0100001011000110: out_v[197] = 10'b1110010011;
    16'b0100001001010110: out_v[197] = 10'b1110011010;
    16'b0110001010000111: out_v[197] = 10'b0101111111;
    16'b0000000000001110: out_v[197] = 10'b0101010100;
    16'b0000000000000101: out_v[197] = 10'b0000110111;
    16'b0100000001010000: out_v[197] = 10'b0111001011;
    16'b0000000001001000: out_v[197] = 10'b0101000100;
    16'b0100000011000010: out_v[197] = 10'b1000100101;
    16'b0110000011000100: out_v[197] = 10'b0110100010;
    16'b0110000011000010: out_v[197] = 10'b0111100000;
    16'b0000001001011110: out_v[197] = 10'b0011001000;
    16'b0000001000001010: out_v[197] = 10'b1111001011;
    16'b0000000010011110: out_v[197] = 10'b1010101011;
    16'b0100001001001110: out_v[197] = 10'b1101100111;
    16'b0000001001001110: out_v[197] = 10'b1011100011;
    16'b0100000001001101: out_v[197] = 10'b1010100101;
    16'b0000000001001110: out_v[197] = 10'b0100111101;
    16'b0100000001001000: out_v[197] = 10'b0100000000;
    16'b0000000001010100: out_v[197] = 10'b0100010110;
    16'b0100000001010110: out_v[197] = 10'b1110011001;
    16'b0000000001011100: out_v[197] = 10'b1111101010;
    16'b0100000001011100: out_v[197] = 10'b0000101110;
    16'b0100001001010100: out_v[197] = 10'b1110000001;
    16'b0110001011010110: out_v[197] = 10'b0111010000;
    default: out_v[197] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000000000000: out_v[198] = 10'b1000110011;
    16'b0001001000001000: out_v[198] = 10'b0111100011;
    16'b0000001000001001: out_v[198] = 10'b0010001101;
    16'b0000000000001000: out_v[198] = 10'b0000000101;
    16'b0000001000001000: out_v[198] = 10'b0110011100;
    16'b0001001000001001: out_v[198] = 10'b0110001011;
    16'b0000001000000000: out_v[198] = 10'b0110011010;
    16'b0001000000001000: out_v[198] = 10'b1101001010;
    16'b0001001000000000: out_v[198] = 10'b0100100001;
    16'b0000000000001001: out_v[198] = 10'b1100010111;
    16'b0001000000000000: out_v[198] = 10'b1100011010;
    16'b0000001000000001: out_v[198] = 10'b0000011111;
    16'b0001001000000001: out_v[198] = 10'b1010001100;
    16'b0000011001001000: out_v[198] = 10'b0111000011;
    16'b0001010001001000: out_v[198] = 10'b0000011111;
    16'b0000010001001000: out_v[198] = 10'b0001100101;
    16'b0000000000000001: out_v[198] = 10'b0101010100;
    16'b0000010001000000: out_v[198] = 10'b1101000000;
    16'b0000010000001000: out_v[198] = 10'b1111110001;
    16'b0001010001000000: out_v[198] = 10'b1100010101;
    16'b0001000000001001: out_v[198] = 10'b1111100000;
    16'b0001011001001000: out_v[198] = 10'b0011110010;
    16'b0001000000100000: out_v[198] = 10'b0010000100;
    16'b0000000000100000: out_v[198] = 10'b0101110110;
    default: out_v[198] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000001100000000: out_v[199] = 10'b1111100110;
    16'b0000001100001000: out_v[199] = 10'b0111001110;
    16'b1000001100001001: out_v[199] = 10'b0001111101;
    16'b1000000000001001: out_v[199] = 10'b0010111011;
    16'b0000000100001000: out_v[199] = 10'b0010001011;
    16'b0000000100001001: out_v[199] = 10'b0100100100;
    16'b0001001101001000: out_v[199] = 10'b0111111001;
    16'b0001001100001001: out_v[199] = 10'b1010011011;
    16'b0000001100001001: out_v[199] = 10'b0011010011;
    16'b0000000000001001: out_v[199] = 10'b0010011001;
    16'b1000001100001000: out_v[199] = 10'b0001010111;
    16'b0001001100001000: out_v[199] = 10'b0000100011;
    16'b0000000000101001: out_v[199] = 10'b1000000001;
    16'b1000000100001001: out_v[199] = 10'b0101000111;
    16'b0000000000001000: out_v[199] = 10'b0011000011;
    16'b1000000100001000: out_v[199] = 10'b1011011011;
    16'b0001000100001001: out_v[199] = 10'b1100101011;
    16'b0000000000000001: out_v[199] = 10'b0101110011;
    16'b0001000000001001: out_v[199] = 10'b1000111110;
    16'b0000001100000001: out_v[199] = 10'b0110100100;
    16'b0001001101001001: out_v[199] = 10'b0001101111;
    16'b1000001101001000: out_v[199] = 10'b1111110110;
    16'b0001001100000000: out_v[199] = 10'b0001100011;
    16'b1000001100000001: out_v[199] = 10'b1101100111;
    16'b1001001101001000: out_v[199] = 10'b1000110011;
    16'b0000000000000000: out_v[199] = 10'b0110010011;
    16'b1000000000001000: out_v[199] = 10'b1010111100;
    16'b0000000100000001: out_v[199] = 10'b1011111111;
    16'b0000000100000000: out_v[199] = 10'b0110100111;
    16'b1000001100000000: out_v[199] = 10'b0110110110;
    16'b1001001100001001: out_v[199] = 10'b1111001011;
    16'b0011001001000000: out_v[199] = 10'b0011010010;
    16'b0011000001000000: out_v[199] = 10'b0011100101;
    16'b0010000001000000: out_v[199] = 10'b0110100111;
    16'b0010001001000000: out_v[199] = 10'b1100110111;
    16'b0011000000000000: out_v[199] = 10'b0101000111;
    16'b0010001101000000: out_v[199] = 10'b1000110110;
    16'b0011001101000000: out_v[199] = 10'b1100001111;
    16'b1011000001000000: out_v[199] = 10'b1111101100;
    16'b1011000000000000: out_v[199] = 10'b1000010111;
    16'b0011001000000000: out_v[199] = 10'b0011010010;
    16'b0011000001100000: out_v[199] = 10'b1011000101;
    16'b0011001001100001: out_v[199] = 10'b1110000100;
    16'b0010000000000000: out_v[199] = 10'b1000011100;
    16'b0011000001000001: out_v[199] = 10'b0110000100;
    16'b0011000001001000: out_v[199] = 10'b1101100101;
    16'b0011001001000001: out_v[199] = 10'b1010001111;
    16'b0011000001100001: out_v[199] = 10'b1110110011;
    16'b0001000001100001: out_v[199] = 10'b1111110010;
    16'b0111000001100001: out_v[199] = 10'b0110110010;
    16'b1011000001001001: out_v[199] = 10'b1100110111;
    16'b1011000001000001: out_v[199] = 10'b1100110101;
    16'b0001000001000000: out_v[199] = 10'b1100010100;
    16'b0001000001000001: out_v[199] = 10'b1101101110;
    16'b1011000001100001: out_v[199] = 10'b0101111011;
    16'b0011000000000001: out_v[199] = 10'b0111000101;
    16'b1011000101000001: out_v[199] = 10'b1111011011;
    16'b1001000001001000: out_v[199] = 10'b1011100110;
    16'b0011001101000001: out_v[199] = 10'b1101100110;
    16'b0010000001000001: out_v[199] = 10'b0001010011;
    16'b0111000001100000: out_v[199] = 10'b1110000111;
    16'b0101000001100001: out_v[199] = 10'b1011110010;
    16'b1011000001001000: out_v[199] = 10'b1011100010;
    16'b0011000001001001: out_v[199] = 10'b0110111010;
    16'b1011000101001001: out_v[199] = 10'b1010100110;
    16'b0010000000000001: out_v[199] = 10'b0000101000;
    16'b0011000000100001: out_v[199] = 10'b1011101011;
    16'b0011000101000000: out_v[199] = 10'b0110001001;
    16'b1001000001001001: out_v[199] = 10'b1001110110;
    16'b0011000101000001: out_v[199] = 10'b0001010100;
    16'b0010000001100001: out_v[199] = 10'b0111010010;
    16'b1000001000000001: out_v[199] = 10'b0011011100;
    16'b0010001000100000: out_v[199] = 10'b1110110101;
    16'b1000001000000000: out_v[199] = 10'b1111011110;
    16'b0110001100100001: out_v[199] = 10'b0100001101;
    16'b0000001000000000: out_v[199] = 10'b1001001101;
    16'b0000001000000001: out_v[199] = 10'b1000101100;
    16'b0000001000100001: out_v[199] = 10'b0001110001;
    16'b1010001000000000: out_v[199] = 10'b1111001111;
    16'b0010001000000000: out_v[199] = 10'b0001011000;
    16'b1010000000000000: out_v[199] = 10'b1101110100;
    16'b0110001000100001: out_v[199] = 10'b1101101001;
    16'b0010001000000001: out_v[199] = 10'b0011011001;
    16'b0010001100000001: out_v[199] = 10'b0010111111;
    16'b0010001100000000: out_v[199] = 10'b0000110100;
    16'b0010001000100001: out_v[199] = 10'b0011111101;
    16'b0110001000000001: out_v[199] = 10'b0101111111;
    16'b0000001000100000: out_v[199] = 10'b1010111100;
    16'b0100001000100001: out_v[199] = 10'b1000110010;
    16'b1110001000100001: out_v[199] = 10'b0011110001;
    16'b0110000000100001: out_v[199] = 10'b0001100011;
    16'b1000000000000000: out_v[199] = 10'b0101101010;
    16'b0100001100100001: out_v[199] = 10'b0010001100;
    16'b1010000000000001: out_v[199] = 10'b0011110100;
    16'b0010000000100001: out_v[199] = 10'b1011110011;
    16'b1000001000100001: out_v[199] = 10'b0000110110;
    16'b0000001100100001: out_v[199] = 10'b0110111110;
    16'b1010000000001000: out_v[199] = 10'b1101001110;
    16'b1100001000100001: out_v[199] = 10'b1111110111;
    16'b0010000000100000: out_v[199] = 10'b1101000110;
    16'b1010001000000001: out_v[199] = 10'b0111111011;
    16'b0000001100100000: out_v[199] = 10'b1011011011;
    16'b0010000101001000: out_v[199] = 10'b0110110110;
    16'b0010001101001000: out_v[199] = 10'b1010101100;
    16'b0010000001001000: out_v[199] = 10'b1011010110;
    16'b0010000101000000: out_v[199] = 10'b0001011101;
    16'b0011001101001000: out_v[199] = 10'b0011011000;
    16'b0010000100000000: out_v[199] = 10'b1000111110;
    16'b0010000000001000: out_v[199] = 10'b1100011110;
    16'b0000000001000000: out_v[199] = 10'b0011110111;
    16'b0011000101001000: out_v[199] = 10'b1101111111;
    16'b0010000100001000: out_v[199] = 10'b1100010010;
    16'b0001001101000000: out_v[199] = 10'b1001110010;
    16'b0010000001100000: out_v[199] = 10'b0010000100;
    16'b0001000001001000: out_v[199] = 10'b1101011110;
    16'b0001000101000000: out_v[199] = 10'b1000111000;
    16'b0000001101000000: out_v[199] = 10'b0011000101;
    16'b1010001101000000: out_v[199] = 10'b0111010001;
    16'b1010000100000000: out_v[199] = 10'b1011011111;
    16'b0010000100000001: out_v[199] = 10'b0001101010;
    16'b0011001001001000: out_v[199] = 10'b0110000010;
    16'b1010001100000000: out_v[199] = 10'b0001111110;
    16'b1010001100000001: out_v[199] = 10'b1111100001;
    16'b0001001000000000: out_v[199] = 10'b1000101000;
    16'b0001001100000001: out_v[199] = 10'b1011101011;
    16'b0001001101000001: out_v[199] = 10'b1001111010;
    16'b0011001100000001: out_v[199] = 10'b1110010101;
    16'b0001000101000001: out_v[199] = 10'b0011111000;
    16'b0011001100000000: out_v[199] = 10'b1100010110;
    16'b0011000101001001: out_v[199] = 10'b1111101110;
    16'b0011000001101001: out_v[199] = 10'b0101100011;
    16'b0011000100000001: out_v[199] = 10'b0010011001;
    16'b0011000000001001: out_v[199] = 10'b0001010111;
    16'b0010000001001001: out_v[199] = 10'b1101000011;
    16'b0011000100000000: out_v[199] = 10'b0100101001;
    16'b0011001101001001: out_v[199] = 10'b1010110011;
    16'b0000000101000000: out_v[199] = 10'b0111011100;
    16'b0000000101001000: out_v[199] = 10'b1001110011;
    16'b0000001101001000: out_v[199] = 10'b1001001011;
    16'b0000000001001000: out_v[199] = 10'b0010010000;
    16'b0110000001000000: out_v[199] = 10'b0111110011;
    16'b0001000101001000: out_v[199] = 10'b1100001110;
    16'b0010001100001000: out_v[199] = 10'b1101000101;
    16'b1011001101001000: out_v[199] = 10'b0101010110;
    16'b0011001000000001: out_v[199] = 10'b0100110101;
    16'b1010001101001000: out_v[199] = 10'b0111110011;
    16'b0010000000001001: out_v[199] = 10'b1110000110;
    16'b0011001100001000: out_v[199] = 10'b0110010111;
    default: out_v[199] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000110101000: out_v[200] = 10'b0011010111;
    16'b0100000110101001: out_v[200] = 10'b0110001111;
    16'b0100000100101101: out_v[200] = 10'b1011000011;
    16'b0100000100001101: out_v[200] = 10'b0000010001;
    16'b0100000110101000: out_v[200] = 10'b0001011111;
    16'b0000000100101101: out_v[200] = 10'b1000000011;
    16'b0000000100001101: out_v[200] = 10'b1001110001;
    16'b0000000000001101: out_v[200] = 10'b1001010011;
    16'b0000000110101001: out_v[200] = 10'b1101010010;
    16'b0100000110101101: out_v[200] = 10'b0001000001;
    16'b0100000110001000: out_v[200] = 10'b0011000001;
    16'b0100000010001000: out_v[200] = 10'b1000011001;
    16'b0100000110001101: out_v[200] = 10'b0100111111;
    16'b0100000110100000: out_v[200] = 10'b0111101011;
    16'b0100000100001001: out_v[200] = 10'b1111100011;
    16'b0100000100000101: out_v[200] = 10'b0100101111;
    16'b0100000000001101: out_v[200] = 10'b0101001011;
    16'b0100000110100101: out_v[200] = 10'b1011001101;
    16'b0100000110100001: out_v[200] = 10'b1010100011;
    16'b0100000010101001: out_v[200] = 10'b0110010011;
    16'b0100000110001001: out_v[200] = 10'b0001101011;
    16'b0100000010100001: out_v[200] = 10'b1111010011;
    16'b0000000000000101: out_v[200] = 10'b0011011011;
    16'b0100000100101001: out_v[200] = 10'b0110110000;
    16'b0100000000000101: out_v[200] = 10'b1101111001;
    16'b0000000110100001: out_v[200] = 10'b1011011110;
    16'b0000000110001000: out_v[200] = 10'b0011100011;
    16'b0100000010101101: out_v[200] = 10'b0010111011;
    16'b0100000000001001: out_v[200] = 10'b1110011011;
    16'b0000000110100000: out_v[200] = 10'b0111100111;
    16'b0000000010001000: out_v[200] = 10'b1100111001;
    16'b0100000100100101: out_v[200] = 10'b0101001011;
    16'b0100000110101100: out_v[200] = 10'b1000101111;
    16'b0000000100101000: out_v[200] = 10'b1000101110;
    16'b0100000010000000: out_v[200] = 10'b0010110011;
    16'b0000000100000101: out_v[200] = 10'b1000011111;
    16'b0000000110101101: out_v[200] = 10'b0110011011;
    16'b0100000110000000: out_v[200] = 10'b0100100011;
    16'b0010000000000000: out_v[200] = 10'b1000011010;
    16'b0010000100000000: out_v[200] = 10'b0010100100;
    16'b0010000100100000: out_v[200] = 10'b1100000000;
    16'b0010000100101000: out_v[200] = 10'b0100110100;
    16'b0010000000100000: out_v[200] = 10'b1111010000;
    16'b0000000000000000: out_v[200] = 10'b1011000100;
    16'b0000000000001000: out_v[200] = 10'b0010001110;
    16'b0010000000001000: out_v[200] = 10'b0110011111;
    16'b0010010000000000: out_v[200] = 10'b1000111100;
    16'b0010000110001001: out_v[200] = 10'b0011000111;
    16'b0000000100000000: out_v[200] = 10'b0110000100;
    16'b0010010000001001: out_v[200] = 10'b1001110110;
    16'b0010000100001000: out_v[200] = 10'b0100011110;
    16'b0000010000001000: out_v[200] = 10'b1010000101;
    16'b0010000110000001: out_v[200] = 10'b0110100110;
    16'b0010000010000001: out_v[200] = 10'b1110000100;
    16'b0000000100001000: out_v[200] = 10'b0110010010;
    16'b0010000010001000: out_v[200] = 10'b0011011100;
    16'b0110010010001001: out_v[200] = 10'b0010111111;
    16'b0000000000001001: out_v[200] = 10'b1100111010;
    16'b0010000110101001: out_v[200] = 10'b0111101110;
    16'b0000010000001001: out_v[200] = 10'b0011111110;
    16'b0010000010001001: out_v[200] = 10'b0011101111;
    16'b0000010010001001: out_v[200] = 10'b0010110101;
    16'b0110000010001001: out_v[200] = 10'b1010100110;
    16'b0010010010000001: out_v[200] = 10'b0111110010;
    16'b0110000010000001: out_v[200] = 10'b0110010100;
    16'b0000000100001001: out_v[200] = 10'b1111110011;
    16'b0000000000000001: out_v[200] = 10'b0010110101;
    16'b0010000000001001: out_v[200] = 10'b0011011001;
    16'b0010010010001001: out_v[200] = 10'b1101100111;
    16'b0010000100001001: out_v[200] = 10'b1010001101;
    16'b0010010000001000: out_v[200] = 10'b0110110101;
    16'b0010000100101001: out_v[200] = 10'b0010101001;
    16'b0010000100000001: out_v[200] = 10'b1011101101;
    16'b0000000100000001: out_v[200] = 10'b1011011110;
    16'b0000000010001001: out_v[200] = 10'b0000111110;
    16'b0010000110001000: out_v[200] = 10'b1100101010;
    16'b0110000110001001: out_v[200] = 10'b1011011110;
    16'b0000000110001001: out_v[200] = 10'b0110010110;
    16'b0010010010001000: out_v[200] = 10'b0011000011;
    16'b0010000000000001: out_v[200] = 10'b0001110001;
    16'b0010000110000000: out_v[200] = 10'b1001101000;
    16'b0110000110000001: out_v[200] = 10'b1111010110;
    16'b0000000000101000: out_v[200] = 10'b0011101100;
    16'b0000000100100000: out_v[200] = 10'b0001101101;
    16'b0100000000101001: out_v[200] = 10'b1011111110;
    16'b0010000110101000: out_v[200] = 10'b1011011000;
    16'b0000000010101000: out_v[200] = 10'b0111000101;
    16'b0100000000101000: out_v[200] = 10'b1011100001;
    16'b0010000000101000: out_v[200] = 10'b1110000011;
    16'b0110000110101000: out_v[200] = 10'b1001011011;
    16'b0100000100101000: out_v[200] = 10'b1010010100;
    16'b0010000010101000: out_v[200] = 10'b1101101110;
    16'b0000000100101001: out_v[200] = 10'b0001100100;
    16'b0000000000100000: out_v[200] = 10'b1011100001;
    16'b0100000100100000: out_v[200] = 10'b1001001010;
    16'b0010000010000000: out_v[200] = 10'b0011111010;
    16'b0000010000101001: out_v[200] = 10'b0111001111;
    16'b0100000010101000: out_v[200] = 10'b1111100110;
    16'b0100000000100000: out_v[200] = 10'b1100100010;
    16'b0000010000101000: out_v[200] = 10'b1111111000;
    16'b0000000000101001: out_v[200] = 10'b0011101110;
    16'b0010000010100001: out_v[200] = 10'b0010011111;
    16'b0010000010100000: out_v[200] = 10'b1000100110;
    16'b0110000010100000: out_v[200] = 10'b1110001110;
    16'b0110000010000000: out_v[200] = 10'b0100111011;
    16'b0010000110100000: out_v[200] = 10'b0001010100;
    16'b0110000110100000: out_v[200] = 10'b0000111100;
    16'b0110000010001000: out_v[200] = 10'b0011111001;
    16'b0000000010000000: out_v[200] = 10'b0100010011;
    16'b0010000010001010: out_v[200] = 10'b1011111111;
    16'b0110000110100001: out_v[200] = 10'b0111110010;
    16'b0000000010100000: out_v[200] = 10'b1100100010;
    16'b0110000110100100: out_v[200] = 10'b0100110010;
    16'b0110000010000100: out_v[200] = 10'b1001011100;
    16'b0110000110000000: out_v[200] = 10'b0111100000;
    16'b0110000010100001: out_v[200] = 10'b1111100010;
    16'b0000000110000000: out_v[200] = 10'b1000110011;
    16'b0010000110100001: out_v[200] = 10'b1100011110;
    16'b0000000100100001: out_v[200] = 10'b1000110110;
    16'b0010000000100001: out_v[200] = 10'b1010011100;
    16'b0000000000100001: out_v[200] = 10'b0001111001;
    16'b0010000100100001: out_v[200] = 10'b1111111011;
    16'b0000000010100001: out_v[200] = 10'b0001001011;
    16'b0110010010001000: out_v[200] = 10'b0001101001;
    16'b0110000010001100: out_v[200] = 10'b1001010110;
    16'b0110000110101101: out_v[200] = 10'b1111010011;
    16'b0110010110101000: out_v[200] = 10'b1110110001;
    16'b0110000110001000: out_v[200] = 10'b1001111010;
    16'b0100010110101000: out_v[200] = 10'b1111110101;
    16'b0100000010001100: out_v[200] = 10'b1111000111;
    16'b0110010110001000: out_v[200] = 10'b1100101111;
    16'b0110010010001100: out_v[200] = 10'b1110011111;
    16'b0110000110101001: out_v[200] = 10'b1101001000;
    16'b0010010100101000: out_v[200] = 10'b1111000011;
    16'b0110000110101100: out_v[200] = 10'b0011011110;
    16'b0110000000001101: out_v[200] = 10'b0011111111;
    16'b0100010010001000: out_v[200] = 10'b1111001110;
    16'b0010010110101000: out_v[200] = 10'b1111110100;
    16'b0110010110101100: out_v[200] = 10'b1001110100;
    16'b0100000100000000: out_v[200] = 10'b0010101011;
    16'b0100000100001000: out_v[200] = 10'b0111100110;
    16'b0110000100000000: out_v[200] = 10'b1011100001;
    16'b0110000100100000: out_v[200] = 10'b1100011111;
    16'b0010000110001010: out_v[200] = 10'b1100111110;
    16'b0000000110001010: out_v[200] = 10'b1101001111;
    default: out_v[200] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000010000001100: out_v[201] = 10'b0100001010;
    16'b0000001000001101: out_v[201] = 10'b0010110101;
    16'b0001001000001101: out_v[201] = 10'b0001100001;
    16'b0001011000001101: out_v[201] = 10'b1110110011;
    16'b0000000000001101: out_v[201] = 10'b0001000101;
    16'b0001000000001101: out_v[201] = 10'b0001100011;
    16'b0000000000000001: out_v[201] = 10'b0000001111;
    16'b0000011000001101: out_v[201] = 10'b0111011110;
    16'b0000010000001101: out_v[201] = 10'b1101001110;
    16'b0000011000001001: out_v[201] = 10'b1111101111;
    16'b0000010000001001: out_v[201] = 10'b0011010101;
    16'b0000010000001000: out_v[201] = 10'b1100000111;
    16'b0000011000001100: out_v[201] = 10'b1001100100;
    16'b0001010000001101: out_v[201] = 10'b0100000011;
    16'b0000011000000101: out_v[201] = 10'b1011011110;
    16'b0000000000000101: out_v[201] = 10'b0110011010;
    16'b0000001000011101: out_v[201] = 10'b1011011101;
    16'b0000001000000101: out_v[201] = 10'b1110000001;
    16'b0000010000000100: out_v[201] = 10'b0000001111;
    16'b0000001000000001: out_v[201] = 10'b0010010001;
    16'b0001010000001001: out_v[201] = 10'b0000011011;
    16'b0000001000010101: out_v[201] = 10'b1011010001;
    16'b0000010000000101: out_v[201] = 10'b1011000100;
    16'b0000000000001001: out_v[201] = 10'b0001010011;
    16'b0000000000001100: out_v[201] = 10'b1100100111;
    16'b0000001000001001: out_v[201] = 10'b1000100101;
    16'b0000011000011101: out_v[201] = 10'b1110111110;
    16'b0001000000001100: out_v[201] = 10'b0100111110;
    16'b0001011000001001: out_v[201] = 10'b0111111101;
    16'b0000000000010100: out_v[201] = 10'b0101011000;
    16'b0000000000000100: out_v[201] = 10'b0011010010;
    16'b0000000000001000: out_v[201] = 10'b1101001110;
    16'b0000000000000000: out_v[201] = 10'b0110010000;
    16'b0000001000010100: out_v[201] = 10'b1110001001;
    16'b0000010000000000: out_v[201] = 10'b1101001011;
    16'b0000000000010000: out_v[201] = 10'b1001011010;
    16'b0000001000010000: out_v[201] = 10'b0111000111;
    16'b0000001000000100: out_v[201] = 10'b0110110000;
    16'b0000001000000000: out_v[201] = 10'b1000000010;
    16'b0000001000001100: out_v[201] = 10'b0010100101;
    16'b0000011000010001: out_v[201] = 10'b1010110101;
    16'b0000010000000001: out_v[201] = 10'b1111001011;
    16'b0000011000000001: out_v[201] = 10'b1111000011;
    16'b0000011000000100: out_v[201] = 10'b1110001011;
    16'b0000011000001000: out_v[201] = 10'b1100000010;
    16'b0000011000011001: out_v[201] = 10'b0000001111;
    16'b0000011000011100: out_v[201] = 10'b0000101101;
    16'b0000011000010101: out_v[201] = 10'b1010111101;
    16'b0000011000000000: out_v[201] = 10'b1111011100;
    16'b0000000010001000: out_v[201] = 10'b1011000001;
    16'b0000111000001100: out_v[201] = 10'b1000010011;
    16'b0000010000000010: out_v[201] = 10'b0100101010;
    16'b0000000010000010: out_v[201] = 10'b0101111111;
    16'b0000000000001110: out_v[201] = 10'b0101111110;
    16'b0000000000000010: out_v[201] = 10'b1000101011;
    16'b0000001000001000: out_v[201] = 10'b0101110011;
    16'b0000000000001010: out_v[201] = 10'b0011110001;
    16'b0000000000001011: out_v[201] = 10'b0110010101;
    16'b0001001000000001: out_v[201] = 10'b1100011110;
    16'b0000000010000000: out_v[201] = 10'b1100001010;
    16'b0001000000001011: out_v[201] = 10'b0101111101;
    16'b0001001000001001: out_v[201] = 10'b1100110111;
    16'b0000000010001001: out_v[201] = 10'b0111010100;
    16'b0001001000000101: out_v[201] = 10'b1101101110;
    16'b0000000000010101: out_v[201] = 10'b1011010000;
    16'b0001000000000001: out_v[201] = 10'b1101010011;
    16'b0000000000000011: out_v[201] = 10'b1000001011;
    16'b0000001000011001: out_v[201] = 10'b1001101101;
    16'b0000001010001000: out_v[201] = 10'b0011110101;
    16'b0001001000001011: out_v[201] = 10'b1011111011;
    16'b0001000000001001: out_v[201] = 10'b0100011011;
    16'b0001000000000011: out_v[201] = 10'b1001111001;
    16'b0000001010001001: out_v[201] = 10'b0111010110;
    16'b0001001000011001: out_v[201] = 10'b0111111111;
    16'b0000000000011100: out_v[201] = 10'b1100100011;
    16'b0000001000011100: out_v[201] = 10'b1100101110;
    16'b0000010000011100: out_v[201] = 10'b1100110000;
    16'b0000010000011101: out_v[201] = 10'b1010100111;
    16'b0000000000100001: out_v[201] = 10'b0111000111;
    16'b0000000000011101: out_v[201] = 10'b1011000010;
    16'b0001000010001000: out_v[201] = 10'b0111010011;
    16'b0001001000001100: out_v[201] = 10'b1111100010;
    16'b0000000010001100: out_v[201] = 10'b0110110010;
    16'b0000000010001010: out_v[201] = 10'b1011101001;
    16'b0000000010000100: out_v[201] = 10'b0101110110;
    16'b0001000000001000: out_v[201] = 10'b0011000010;
    16'b0100000000000100: out_v[201] = 10'b1100001011;
    16'b0001000000000100: out_v[201] = 10'b1110000111;
    16'b0001001000000100: out_v[201] = 10'b1011101111;
    16'b0000010000001110: out_v[201] = 10'b1000110111;
    16'b0000010000000110: out_v[201] = 10'b1010011111;
    16'b0000000000000110: out_v[201] = 10'b0101100111;
    16'b0000000010001011: out_v[201] = 10'b1111100011;
    16'b1001000000000001: out_v[201] = 10'b1011000000;
    16'b0001000010001001: out_v[201] = 10'b1001110110;
    default: out_v[201] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000011000100100: out_v[202] = 10'b0111110011;
    16'b1000011000100100: out_v[202] = 10'b1010100011;
    16'b1100011000100110: out_v[202] = 10'b0101101011;
    16'b0000001000100100: out_v[202] = 10'b0111000011;
    16'b0000010000100100: out_v[202] = 10'b1001010001;
    16'b0100010000010110: out_v[202] = 10'b1011001001;
    16'b1000010000100100: out_v[202] = 10'b1001100001;
    16'b0000010000100000: out_v[202] = 10'b1100100101;
    16'b1000000000000100: out_v[202] = 10'b1010011010;
    16'b0100001000100100: out_v[202] = 10'b0110100011;
    16'b0000010000000100: out_v[202] = 10'b0011101011;
    16'b1000011000100000: out_v[202] = 10'b0111110011;
    16'b0000011000100000: out_v[202] = 10'b1101110010;
    16'b0000001000000100: out_v[202] = 10'b0110000001;
    16'b1000001000100100: out_v[202] = 10'b0010011101;
    16'b1000000000100100: out_v[202] = 10'b1100010100;
    16'b0100001000000110: out_v[202] = 10'b1000011110;
    16'b1000010000000100: out_v[202] = 10'b1100001000;
    16'b0100001000010110: out_v[202] = 10'b0010101010;
    16'b0100000000000110: out_v[202] = 10'b1011100011;
    16'b0100001000000100: out_v[202] = 10'b1000110111;
    16'b0000000000100100: out_v[202] = 10'b1001011011;
    16'b0100000000010110: out_v[202] = 10'b1001101111;
    16'b1000010000100000: out_v[202] = 10'b0100110001;
    16'b0000000000000100: out_v[202] = 10'b1001111010;
    16'b0100010000000110: out_v[202] = 10'b0101110101;
    16'b0100011000100110: out_v[202] = 10'b1100100011;
    16'b0100011000100100: out_v[202] = 10'b0100011001;
    16'b1000001000100000: out_v[202] = 10'b1011101001;
    16'b1100001000000110: out_v[202] = 10'b0110011111;
    16'b0000001000100000: out_v[202] = 10'b0010011100;
    16'b0100001000100110: out_v[202] = 10'b0110100011;
    16'b0100011000110110: out_v[202] = 10'b0101100001;
    16'b1100011000000110: out_v[202] = 10'b0111011011;
    16'b1000011000000000: out_v[202] = 10'b0101011111;
    16'b0100011000010110: out_v[202] = 10'b0000110111;
    16'b1100011000100100: out_v[202] = 10'b0001111101;
    16'b1100001000010110: out_v[202] = 10'b1011111011;
    16'b0000011000000100: out_v[202] = 10'b1110111010;
    16'b0000011000000000: out_v[202] = 10'b0100110110;
    16'b0000010000000000: out_v[202] = 10'b1101011101;
    16'b1000000000000000: out_v[202] = 10'b1010001111;
    16'b0000000000000000: out_v[202] = 10'b1001111011;
    16'b1000010000010100: out_v[202] = 10'b0111110011;
    16'b1000000000110100: out_v[202] = 10'b1000100110;
    16'b1100000000010100: out_v[202] = 10'b0011100101;
    16'b0000000000100000: out_v[202] = 10'b0000110010;
    16'b1000000000010100: out_v[202] = 10'b0100010101;
    16'b0000000000010100: out_v[202] = 10'b1011011010;
    16'b0100010000010010: out_v[202] = 10'b0100101011;
    16'b0100000000010000: out_v[202] = 10'b0100100111;
    16'b1100000000000100: out_v[202] = 10'b1011110011;
    16'b1100000000100100: out_v[202] = 10'b1001011110;
    16'b0100000000000000: out_v[202] = 10'b1000010011;
    16'b0000010000110000: out_v[202] = 10'b0100010001;
    16'b0000000000001000: out_v[202] = 10'b0100110101;
    16'b0000000000010000: out_v[202] = 10'b1000101100;
    16'b0100000000110000: out_v[202] = 10'b0011011110;
    16'b0100000000000100: out_v[202] = 10'b1101100100;
    16'b0000010000010000: out_v[202] = 10'b0001001101;
    16'b0000000000110000: out_v[202] = 10'b0111001001;
    16'b1100010000000100: out_v[202] = 10'b1001011111;
    16'b1100000000010110: out_v[202] = 10'b0010101110;
    16'b0000010000010100: out_v[202] = 10'b1100001100;
    16'b1000010000000000: out_v[202] = 10'b0011001101;
    16'b1000000000010000: out_v[202] = 10'b0101011110;
    16'b1000001000000100: out_v[202] = 10'b1001010111;
    16'b0100010000000100: out_v[202] = 10'b1010110000;
    16'b1100001000000100: out_v[202] = 10'b1001011101;
    16'b0100010000010100: out_v[202] = 10'b1001011101;
    16'b0100000000010100: out_v[202] = 10'b1111100010;
    16'b0100010000010000: out_v[202] = 10'b1100111000;
    16'b0000010000110100: out_v[202] = 10'b1001000100;
    16'b1100000000000110: out_v[202] = 10'b0001010111;
    16'b0100010000000000: out_v[202] = 10'b1101011101;
    16'b0000000000110100: out_v[202] = 10'b1111010101;
    16'b1100000000110100: out_v[202] = 10'b1111011110;
    16'b0100000000100100: out_v[202] = 10'b0111010110;
    16'b1000000000001100: out_v[202] = 10'b0110000111;
    16'b0000001000000000: out_v[202] = 10'b1001100101;
    16'b1100001000000000: out_v[202] = 10'b0100110001;
    16'b1100001000000010: out_v[202] = 10'b0010101010;
    16'b0100011000000010: out_v[202] = 10'b0100101000;
    16'b0100011000000100: out_v[202] = 10'b0111101100;
    16'b0100001000000000: out_v[202] = 10'b0110011001;
    16'b0100001000000010: out_v[202] = 10'b0011101011;
    16'b1000001000000000: out_v[202] = 10'b1000100110;
    16'b0100011000100000: out_v[202] = 10'b0110101001;
    16'b1000010000001100: out_v[202] = 10'b1001111000;
    16'b1100011000000000: out_v[202] = 10'b1000011101;
    16'b1100001000100000: out_v[202] = 10'b0001101010;
    16'b1000000000101100: out_v[202] = 10'b1111101101;
    16'b1100001000100100: out_v[202] = 10'b0110111010;
    16'b1000011000000100: out_v[202] = 10'b0011110110;
    16'b0100011000000000: out_v[202] = 10'b0010001100;
    16'b1000000000100000: out_v[202] = 10'b0000111010;
    16'b1100011000100000: out_v[202] = 10'b1110001000;
    16'b1100011000000100: out_v[202] = 10'b1101010110;
    16'b0100001000100000: out_v[202] = 10'b1000001110;
    16'b0100000000100000: out_v[202] = 10'b0011011100;
    16'b0100000000000010: out_v[202] = 10'b1111100001;
    16'b0000000000000010: out_v[202] = 10'b0111101000;
    16'b0100000000100010: out_v[202] = 10'b1001001010;
    16'b0100001000100010: out_v[202] = 10'b1100011001;
    16'b0000000000100010: out_v[202] = 10'b0011010011;
    16'b0100001000110110: out_v[202] = 10'b1110110010;
    16'b0010000000100100: out_v[202] = 10'b1111100100;
    16'b0100000000110010: out_v[202] = 10'b1101110011;
    16'b0010000000000000: out_v[202] = 10'b1001001101;
    16'b0010000000100000: out_v[202] = 10'b0100110111;
    16'b0110000000100100: out_v[202] = 10'b1010101101;
    16'b0010010000100100: out_v[202] = 10'b0111010111;
    16'b0110000000100000: out_v[202] = 10'b1111111111;
    16'b0100000000100110: out_v[202] = 10'b1000111100;
    16'b0000011000000010: out_v[202] = 10'b0011100100;
    16'b0000010000000010: out_v[202] = 10'b1110101100;
    16'b0100010000000011: out_v[202] = 10'b0101100010;
    16'b0100011000000011: out_v[202] = 10'b0110011010;
    16'b0000010000000110: out_v[202] = 10'b0011100101;
    16'b0100011000000001: out_v[202] = 10'b0011101111;
    16'b0100010000000010: out_v[202] = 10'b0010001001;
    16'b0000010000000011: out_v[202] = 10'b0011111111;
    16'b0100011000100010: out_v[202] = 10'b1111000110;
    16'b0100011000000110: out_v[202] = 10'b0011011100;
    16'b1100010000000110: out_v[202] = 10'b0110000101;
    16'b0100010000100000: out_v[202] = 10'b1110000110;
    16'b0100010000000001: out_v[202] = 10'b1001111001;
    16'b0000011000100001: out_v[202] = 10'b0101101011;
    16'b0100010000100010: out_v[202] = 10'b1110100011;
    16'b0000000000100001: out_v[202] = 10'b1010000111;
    16'b0000010000100001: out_v[202] = 10'b1101001011;
    default: out_v[202] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000010000001: out_v[203] = 10'b1001010101;
    16'b1100000000100000: out_v[203] = 10'b1100100010;
    16'b1100000000101001: out_v[203] = 10'b1011010111;
    16'b0000000000101000: out_v[203] = 10'b1010010111;
    16'b0000000000000001: out_v[203] = 10'b1111000000;
    16'b0000000000101001: out_v[203] = 10'b1010011100;
    16'b1100000000100001: out_v[203] = 10'b1101111010;
    16'b0000000000001001: out_v[203] = 10'b0001000100;
    16'b0100000000101000: out_v[203] = 10'b1111010010;
    16'b0100000010101001: out_v[203] = 10'b0001010111;
    16'b0000000010100001: out_v[203] = 10'b0000110111;
    16'b1000000000101000: out_v[203] = 10'b1110001000;
    16'b1000000000100001: out_v[203] = 10'b0011011111;
    16'b0000000010001001: out_v[203] = 10'b1110011010;
    16'b0100000010001000: out_v[203] = 10'b0010111011;
    16'b0000000010101000: out_v[203] = 10'b0110111011;
    16'b0100000000100000: out_v[203] = 10'b1011011111;
    16'b1000000000100000: out_v[203] = 10'b0010010010;
    16'b0000000000100001: out_v[203] = 10'b0111100100;
    16'b0000000010101001: out_v[203] = 10'b0011001011;
    16'b0000000000100000: out_v[203] = 10'b1010110011;
    16'b1000000000001001: out_v[203] = 10'b1000000111;
    16'b0100000000101001: out_v[203] = 10'b0111010101;
    16'b1100000000000001: out_v[203] = 10'b0100100011;
    16'b0000000010000000: out_v[203] = 10'b1000001011;
    16'b1100000000101000: out_v[203] = 10'b1010111111;
    16'b0100000000001000: out_v[203] = 10'b1010111010;
    16'b0000000010001000: out_v[203] = 10'b1010101000;
    16'b0100000010101000: out_v[203] = 10'b0011110010;
    16'b1000000000000001: out_v[203] = 10'b0100110101;
    16'b1000000000101001: out_v[203] = 10'b0101000010;
    16'b0000000000000000: out_v[203] = 10'b1100110101;
    16'b1000000010001000: out_v[203] = 10'b0110001000;
    16'b0100000000000001: out_v[203] = 10'b0100010111;
    16'b0100000000100001: out_v[203] = 10'b0100001000;
    16'b1000000010101001: out_v[203] = 10'b1011101011;
    16'b0000000000001000: out_v[203] = 10'b0011111001;
    16'b1000000010000000: out_v[203] = 10'b1010111011;
    16'b1000000000000000: out_v[203] = 10'b1110011101;
    16'b1000000010100000: out_v[203] = 10'b0010011100;
    16'b1000000010100001: out_v[203] = 10'b1001111101;
    16'b0000000000001011: out_v[203] = 10'b0110110110;
    16'b0000000000000011: out_v[203] = 10'b1001000011;
    16'b0000000010100000: out_v[203] = 10'b0101100110;
    16'b1000000010000001: out_v[203] = 10'b1110010110;
    16'b0000000000100011: out_v[203] = 10'b1110101011;
    16'b1000000000001000: out_v[203] = 10'b1100001101;
    16'b0100000000001001: out_v[203] = 10'b1110110110;
    16'b1000000010101000: out_v[203] = 10'b0110001000;
    16'b1000000010001001: out_v[203] = 10'b0110110010;
    16'b0100000000000000: out_v[203] = 10'b0100111111;
    16'b0100000010000000: out_v[203] = 10'b0001111001;
    16'b1100000010000000: out_v[203] = 10'b0110001111;
    16'b1100000000000000: out_v[203] = 10'b0111110001;
    16'b0000000000101011: out_v[203] = 10'b1111010110;
    16'b1000000000101011: out_v[203] = 10'b0101100000;
    16'b1000000000100011: out_v[203] = 10'b0101110000;
    16'b1000000000000011: out_v[203] = 10'b1011001010;
    16'b1000000000001011: out_v[203] = 10'b1011010010;
    16'b0100000010000001: out_v[203] = 10'b1100110111;
    16'b0100000010100001: out_v[203] = 10'b0101010110;
    16'b1100000010000001: out_v[203] = 10'b1100011101;
    default: out_v[203] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100000010000000: out_v[204] = 10'b0011100111;
    16'b0100000011000000: out_v[204] = 10'b1001100011;
    16'b0100000011001000: out_v[204] = 10'b0101100001;
    16'b0100000010001000: out_v[204] = 10'b1000001101;
    16'b0000000000000000: out_v[204] = 10'b1000000111;
    16'b0100000000000000: out_v[204] = 10'b0011011100;
    16'b0000000001000000: out_v[204] = 10'b1010110011;
    16'b0100000001000000: out_v[204] = 10'b1000110110;
    16'b0000000010000000: out_v[204] = 10'b1100110011;
    16'b0100000000001000: out_v[204] = 10'b1011110010;
    16'b0000000010001000: out_v[204] = 10'b0110100000;
    16'b0000000011000000: out_v[204] = 10'b0101010000;
    16'b0000000000001000: out_v[204] = 10'b1011111100;
    16'b1100000000001100: out_v[204] = 10'b0101010011;
    16'b1000000000001000: out_v[204] = 10'b1110101001;
    16'b0100000000001100: out_v[204] = 10'b0100001011;
    16'b1100000010001000: out_v[204] = 10'b0010000110;
    16'b0100000000000100: out_v[204] = 10'b0001101000;
    16'b1000000010001000: out_v[204] = 10'b0100001101;
    16'b0100000010001100: out_v[204] = 10'b1000011110;
    16'b1100000000001000: out_v[204] = 10'b0011001100;
    16'b1100000000000000: out_v[204] = 10'b1001010111;
    16'b0000000000001100: out_v[204] = 10'b1000001101;
    16'b0101000010001000: out_v[204] = 10'b1000111110;
    16'b0000000011001000: out_v[204] = 10'b0110001011;
    16'b0000000001001000: out_v[204] = 10'b1100110010;
    16'b0100000001001000: out_v[204] = 10'b1010110001;
    16'b0100000100000000: out_v[204] = 10'b0001000000;
    16'b0100100000001000: out_v[204] = 10'b1111000001;
    16'b0000000100000000: out_v[204] = 10'b1101001010;
    16'b0101000000000000: out_v[204] = 10'b0010011001;
    16'b0000000010010000: out_v[204] = 10'b1110000010;
    16'b0001000000000000: out_v[204] = 10'b1110011110;
    16'b0001000010000000: out_v[204] = 10'b0111000000;
    16'b0101000010000000: out_v[204] = 10'b1011001111;
    default: out_v[204] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1000000000100000: out_v[205] = 10'b1011001001;
    16'b1000000000000000: out_v[205] = 10'b1000101111;
    16'b0000000000110100: out_v[205] = 10'b1000110111;
    16'b0000000000100000: out_v[205] = 10'b0100100101;
    16'b0000000000100100: out_v[205] = 10'b1000100111;
    16'b0000000000000100: out_v[205] = 10'b0001000100;
    16'b1000000000110000: out_v[205] = 10'b1011000000;
    16'b0000000000010100: out_v[205] = 10'b0001000010;
    16'b1000000000110100: out_v[205] = 10'b0100100011;
    16'b1000000000100100: out_v[205] = 10'b1111000100;
    16'b1000100000100000: out_v[205] = 10'b1001001011;
    16'b0000000000000000: out_v[205] = 10'b0100010110;
    16'b0000100000100000: out_v[205] = 10'b0101010111;
    16'b0000000000110000: out_v[205] = 10'b1101000000;
    16'b0000100000100100: out_v[205] = 10'b1010100010;
    16'b0000000000010000: out_v[205] = 10'b0101010010;
    16'b1000000000000100: out_v[205] = 10'b1110100111;
    16'b0000100000010000: out_v[205] = 10'b0011010010;
    16'b1000000000010000: out_v[205] = 10'b0110110001;
    16'b0000100000110100: out_v[205] = 10'b0001011100;
    16'b0000100000010100: out_v[205] = 10'b1101001110;
    16'b1000000000010100: out_v[205] = 10'b0000011100;
    16'b1000001010110000: out_v[205] = 10'b1101011000;
    16'b1000001000110000: out_v[205] = 10'b1001000010;
    16'b1000000010110000: out_v[205] = 10'b0101011110;
    16'b0000100000110000: out_v[205] = 10'b0111001000;
    16'b1000000010100000: out_v[205] = 10'b0011111111;
    16'b1000100000110000: out_v[205] = 10'b0001101001;
    16'b1000100000010000: out_v[205] = 10'b1000001011;
    16'b1000001000100000: out_v[205] = 10'b1011011000;
    16'b0000000010110100: out_v[205] = 10'b1111000001;
    16'b0000000010010100: out_v[205] = 10'b0010010001;
    16'b1000001000010000: out_v[205] = 10'b0110011111;
    16'b1000001000010100: out_v[205] = 10'b0000011101;
    16'b1000001010100000: out_v[205] = 10'b0010100011;
    16'b0000001010110100: out_v[205] = 10'b0110011101;
    16'b1000001000110100: out_v[205] = 10'b0111001000;
    16'b0000000010100100: out_v[205] = 10'b1000001100;
    16'b1000000010110100: out_v[205] = 10'b1010111011;
    16'b1000001010010100: out_v[205] = 10'b0001101101;
    16'b1000001010110100: out_v[205] = 10'b0111001001;
    16'b0000000010000100: out_v[205] = 10'b1010100011;
    16'b0000001000110100: out_v[205] = 10'b0011110101;
    16'b1000001000000000: out_v[205] = 10'b1010001010;
    16'b0000000010010000: out_v[205] = 10'b0111001011;
    16'b0000000010000000: out_v[205] = 10'b1101111110;
    16'b0000000010110000: out_v[205] = 10'b1001011110;
    16'b0000001000110000: out_v[205] = 10'b0101101010;
    default: out_v[205] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100000000000001: out_v[206] = 10'b1010010011;
    16'b0000010000000001: out_v[206] = 10'b1001011101;
    16'b0100010100000001: out_v[206] = 10'b1001101101;
    16'b0100000000000000: out_v[206] = 10'b0011110011;
    16'b0100010000000001: out_v[206] = 10'b0100101000;
    16'b0100010000000000: out_v[206] = 10'b0100100101;
    16'b0010010000000001: out_v[206] = 10'b0101000111;
    16'b0110010100000000: out_v[206] = 10'b1111001010;
    16'b0110000000000001: out_v[206] = 10'b0010000011;
    16'b0010010000000000: out_v[206] = 10'b0111100001;
    16'b0000010100000000: out_v[206] = 10'b0100100111;
    16'b0110010000000001: out_v[206] = 10'b0010011011;
    16'b0100010100000000: out_v[206] = 10'b1110110110;
    16'b0000010000001001: out_v[206] = 10'b0001010101;
    16'b0000000000000001: out_v[206] = 10'b1010000001;
    16'b0000010100000001: out_v[206] = 10'b0110011100;
    16'b0110010000000000: out_v[206] = 10'b0010111011;
    16'b0110010100000001: out_v[206] = 10'b1000101011;
    16'b0000010000000000: out_v[206] = 10'b0100101010;
    16'b0000000000000000: out_v[206] = 10'b1000111110;
    16'b0000010100001000: out_v[206] = 10'b0101110000;
    16'b0000000000001001: out_v[206] = 10'b0110010010;
    16'b0100010100001000: out_v[206] = 10'b0101010100;
    16'b0100000000001001: out_v[206] = 10'b1011010010;
    16'b0100010000001001: out_v[206] = 10'b1010101101;
    16'b0000010100001001: out_v[206] = 10'b0010000111;
    16'b0100010100001001: out_v[206] = 10'b1100100110;
    16'b0000000000001000: out_v[206] = 10'b1101011001;
    16'b0100000000001000: out_v[206] = 10'b1100111010;
    16'b0001000000001000: out_v[206] = 10'b0101100100;
    16'b0001010000001001: out_v[206] = 10'b0001000110;
    16'b0000010000001000: out_v[206] = 10'b1100101011;
    16'b0001010000001000: out_v[206] = 10'b0110000101;
    16'b0001010100001001: out_v[206] = 10'b1111110101;
    16'b0100010000001000: out_v[206] = 10'b0101010010;
    16'b0000000100001000: out_v[206] = 10'b1011100110;
    16'b0001000000000000: out_v[206] = 10'b1111000101;
    16'b0001000000001001: out_v[206] = 10'b1001101010;
    16'b0001010000000001: out_v[206] = 10'b0010110111;
    16'b0001010000000000: out_v[206] = 10'b1110101111;
    16'b0001010100001000: out_v[206] = 10'b0111011111;
    16'b0000000100000001: out_v[206] = 10'b1001101101;
    16'b0000000100000000: out_v[206] = 10'b0100001111;
    16'b0000001000001001: out_v[206] = 10'b0110010110;
    16'b0000001000001000: out_v[206] = 10'b0110011111;
    16'b0000000100001001: out_v[206] = 10'b1100101010;
    16'b0000001000000000: out_v[206] = 10'b1101101110;
    16'b0100000100000001: out_v[206] = 10'b0001111111;
    16'b0100001000001001: out_v[206] = 10'b1011001110;
    16'b0000001000000001: out_v[206] = 10'b1110101000;
    16'b0100001000001000: out_v[206] = 10'b1011001000;
    16'b0100000100000000: out_v[206] = 10'b0101110001;
    16'b0100000000001010: out_v[206] = 10'b1111100010;
    16'b0011000000001000: out_v[206] = 10'b1011010111;
    16'b0000000000001010: out_v[206] = 10'b1111111011;
    16'b0101000000000000: out_v[206] = 10'b1011101010;
    16'b0110010000001000: out_v[206] = 10'b0001011110;
    16'b0101000000001000: out_v[206] = 10'b1011000011;
    16'b0100000000000010: out_v[206] = 10'b0111101001;
    16'b0100010000001010: out_v[206] = 10'b1011111011;
    16'b0000000000000010: out_v[206] = 10'b0101010000;
    16'b0010000000001000: out_v[206] = 10'b1101101100;
    16'b0100001000000001: out_v[206] = 10'b0011100110;
    16'b0100001000000000: out_v[206] = 10'b1010001010;
    default: out_v[206] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0011000000000000: out_v[207] = 10'b0010111110;
    16'b0011000000010000: out_v[207] = 10'b1010001011;
    16'b0010010000100000: out_v[207] = 10'b1111000100;
    16'b0110010011100001: out_v[207] = 10'b1110110001;
    16'b0001000001010101: out_v[207] = 10'b0110111110;
    16'b0010010000000001: out_v[207] = 10'b1100100111;
    16'b0010010001100000: out_v[207] = 10'b0010100001;
    16'b0010010001100001: out_v[207] = 10'b0011011111;
    16'b0010000001100001: out_v[207] = 10'b1010000011;
    16'b0010000000000000: out_v[207] = 10'b0111110010;
    16'b0001000000010000: out_v[207] = 10'b0100111001;
    16'b0001010000010000: out_v[207] = 10'b1101000111;
    16'b0110010001100000: out_v[207] = 10'b1101001110;
    16'b0010000000100000: out_v[207] = 10'b0111000101;
    16'b0011000000100000: out_v[207] = 10'b1101100101;
    16'b0011000000100001: out_v[207] = 10'b1010100001;
    16'b0011010000110000: out_v[207] = 10'b1101011000;
    16'b0001100000010100: out_v[207] = 10'b0111100010;
    16'b0001000001010100: out_v[207] = 10'b1000110111;
    16'b0010010000000000: out_v[207] = 10'b1111000000;
    16'b0010010011100001: out_v[207] = 10'b1000111111;
    16'b0001100001010100: out_v[207] = 10'b0001011101;
    16'b0011010000100000: out_v[207] = 10'b0010001011;
    16'b0110010001100001: out_v[207] = 10'b1000111111;
    16'b0001100001010101: out_v[207] = 10'b1111010011;
    16'b0011000000110000: out_v[207] = 10'b0101101111;
    16'b0110010010100001: out_v[207] = 10'b0000011011;
    16'b0010010010100001: out_v[207] = 10'b1011100011;
    16'b0010010000100001: out_v[207] = 10'b1000100110;
    16'b0011000001010001: out_v[207] = 10'b0111111101;
    16'b0011000001110000: out_v[207] = 10'b0011001110;
    16'b0011010000000000: out_v[207] = 10'b0110010001;
    16'b0001000000010100: out_v[207] = 10'b0110100011;
    16'b0001100001110100: out_v[207] = 10'b0010111111;
    16'b0001100000010000: out_v[207] = 10'b1101001010;
    16'b0001000000000000: out_v[207] = 10'b0011011001;
    16'b0011000001110001: out_v[207] = 10'b1111101010;
    16'b0000000000000000: out_v[207] = 10'b1100001111;
    16'b0011010000010000: out_v[207] = 10'b1001011010;
    16'b0001100000110100: out_v[207] = 10'b1011110011;
    16'b0000010000000000: out_v[207] = 10'b1000000011;
    16'b0000010000100000: out_v[207] = 10'b1001001011;
    16'b0001010000100000: out_v[207] = 10'b1010110110;
    16'b0001010000000000: out_v[207] = 10'b0100101101;
    16'b0000010010000000: out_v[207] = 10'b1010110011;
    16'b0000010010000001: out_v[207] = 10'b0000011110;
    16'b0000010000000001: out_v[207] = 10'b1111100100;
    16'b0000000010000001: out_v[207] = 10'b1001111010;
    16'b0001000000100000: out_v[207] = 10'b0101011111;
    16'b0011010000100100: out_v[207] = 10'b0000100111;
    16'b0011010000110100: out_v[207] = 10'b1110100101;
    16'b0001010000110100: out_v[207] = 10'b0110010101;
    16'b0001110000110100: out_v[207] = 10'b1101010011;
    16'b0001010000100100: out_v[207] = 10'b0110001000;
    16'b0011000000100100: out_v[207] = 10'b1100000011;
    16'b0010110000110100: out_v[207] = 10'b1101100101;
    16'b0011100000010000: out_v[207] = 10'b1110001111;
    16'b0001010000000100: out_v[207] = 10'b0101011100;
    16'b0011000000110100: out_v[207] = 10'b1011110111;
    16'b0011110000110100: out_v[207] = 10'b1000101011;
    16'b0011000000010100: out_v[207] = 10'b0011111100;
    16'b0011100000100000: out_v[207] = 10'b1000100111;
    16'b0010010000010000: out_v[207] = 10'b0000001110;
    16'b0011100000110000: out_v[207] = 10'b0111000100;
    16'b0011010000000100: out_v[207] = 10'b1010001100;
    16'b0011100000110100: out_v[207] = 10'b1000010101;
    16'b0011100000010100: out_v[207] = 10'b0111101011;
    16'b0001000000100100: out_v[207] = 10'b1111001001;
    16'b0011000000000100: out_v[207] = 10'b0001100110;
    16'b0010110000010000: out_v[207] = 10'b0010000010;
    16'b0011010000010100: out_v[207] = 10'b1111000001;
    16'b0001000000110100: out_v[207] = 10'b1011001001;
    16'b0011110000110000: out_v[207] = 10'b1001011101;
    16'b0001100000110000: out_v[207] = 10'b1001111111;
    16'b0011110000010100: out_v[207] = 10'b1010100101;
    16'b0010110000110000: out_v[207] = 10'b0010010000;
    16'b0001000000110000: out_v[207] = 10'b1010100111;
    16'b0011110000010000: out_v[207] = 10'b1111001010;
    16'b0001000000000100: out_v[207] = 10'b0011001111;
    16'b0001110000010000: out_v[207] = 10'b1001100011;
    16'b0010000000010000: out_v[207] = 10'b0101010010;
    16'b0001110000000100: out_v[207] = 10'b1100001000;
    16'b0000110000010100: out_v[207] = 10'b1111101000;
    16'b0001110000010100: out_v[207] = 10'b1111010100;
    16'b0001110000000000: out_v[207] = 10'b0001110110;
    16'b0111010000100000: out_v[207] = 10'b1100001011;
    16'b0000110000010000: out_v[207] = 10'b0010110000;
    16'b0010100000010000: out_v[207] = 10'b0110001111;
    16'b0011110000000000: out_v[207] = 10'b0011110001;
    16'b0010000000100001: out_v[207] = 10'b1010110011;
    16'b0000000010100000: out_v[207] = 10'b0101111100;
    16'b0010000010100001: out_v[207] = 10'b0110011000;
    16'b0000000000100000: out_v[207] = 10'b1111000101;
    16'b0010100000010001: out_v[207] = 10'b0101011011;
    16'b0000000000010000: out_v[207] = 10'b0100110110;
    16'b0010100000000000: out_v[207] = 10'b0110000010;
    16'b0010000000110001: out_v[207] = 10'b0101010110;
    16'b0000000000100001: out_v[207] = 10'b0001011010;
    16'b0000000010100001: out_v[207] = 10'b0110100110;
    16'b0000000000110000: out_v[207] = 10'b1111000111;
    16'b0000000000000001: out_v[207] = 10'b0011110010;
    16'b0010110000000000: out_v[207] = 10'b0001110011;
    16'b0010000000110000: out_v[207] = 10'b1101011011;
    16'b0000010000110000: out_v[207] = 10'b0011110001;
    16'b0010000000000001: out_v[207] = 10'b0111010011;
    16'b0010000000010001: out_v[207] = 10'b0100111010;
    16'b0010100010010001: out_v[207] = 10'b1111001111;
    16'b0010000010010001: out_v[207] = 10'b1100011010;
    16'b0000010000010000: out_v[207] = 10'b1001001101;
    16'b0010000010110001: out_v[207] = 10'b1100100100;
    16'b0010000010000001: out_v[207] = 10'b0110010111;
    16'b0000010001100000: out_v[207] = 10'b1100110010;
    16'b0010010010000001: out_v[207] = 10'b1001000111;
    16'b0000010010100001: out_v[207] = 10'b0101100100;
    16'b0000010000100001: out_v[207] = 10'b0001100100;
    16'b0011000000000001: out_v[207] = 10'b1011111110;
    16'b0000010001000000: out_v[207] = 10'b0111100100;
    16'b0010000010000000: out_v[207] = 10'b0011101010;
    16'b0000100000010100: out_v[207] = 10'b0000111111;
    16'b0011000010000000: out_v[207] = 10'b0100110111;
    16'b0011000010010001: out_v[207] = 10'b0111011001;
    16'b0011000010000001: out_v[207] = 10'b0011001110;
    16'b0010010000010001: out_v[207] = 10'b0100100111;
    16'b0011000000010001: out_v[207] = 10'b0000001111;
    16'b0010100000110000: out_v[207] = 10'b1111001011;
    16'b0011000001100000: out_v[207] = 10'b1001110000;
    16'b0010100001110000: out_v[207] = 10'b1001101010;
    16'b0010010010100000: out_v[207] = 10'b1100100010;
    16'b0000100000110000: out_v[207] = 10'b0100100111;
    16'b0010010000110000: out_v[207] = 10'b1100001101;
    16'b1000010000110000: out_v[207] = 10'b1100101101;
    16'b0000110000110000: out_v[207] = 10'b0011110100;
    16'b1000010000100001: out_v[207] = 10'b0111001001;
    16'b1000010000100000: out_v[207] = 10'b0101000111;
    16'b1010110000110000: out_v[207] = 10'b0111101101;
    16'b1000110000110000: out_v[207] = 10'b1100010011;
    16'b0010011000000000: out_v[207] = 10'b1001000111;
    16'b0000100000010000: out_v[207] = 10'b1000101011;
    16'b0010111000010000: out_v[207] = 10'b0000111110;
    16'b0010110000110001: out_v[207] = 10'b1011011010;
    16'b1000000000110000: out_v[207] = 10'b1100111110;
    16'b0010010000110001: out_v[207] = 10'b0010111100;
    16'b0001000000100001: out_v[207] = 10'b0010101111;
    16'b0011100000010001: out_v[207] = 10'b1101100001;
    16'b0011010000010001: out_v[207] = 10'b0110010011;
    16'b0001000000000001: out_v[207] = 10'b1011010101;
    16'b1000000000100000: out_v[207] = 10'b1101111111;
    default: out_v[207] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001000000001100: out_v[208] = 10'b1101010110;
    16'b0000000010011100: out_v[208] = 10'b0111110111;
    16'b0001000010011000: out_v[208] = 10'b1101001011;
    16'b0001000000011000: out_v[208] = 10'b1100100011;
    16'b0001010000011000: out_v[208] = 10'b1011101001;
    16'b0001000010011100: out_v[208] = 10'b0101001111;
    16'b0001010000000000: out_v[208] = 10'b0101010011;
    16'b0001010010001000: out_v[208] = 10'b1110010111;
    16'b0000000000001000: out_v[208] = 10'b0001010111;
    16'b0001000000001000: out_v[208] = 10'b1011101111;
    16'b0001010010011000: out_v[208] = 10'b1000110100;
    16'b0000000000011100: out_v[208] = 10'b1100000111;
    16'b0001000000011100: out_v[208] = 10'b1101001010;
    16'b0000000000011000: out_v[208] = 10'b0110111000;
    16'b0000010000011000: out_v[208] = 10'b0100110011;
    16'b0001010000001000: out_v[208] = 10'b1110101111;
    16'b0000000010010100: out_v[208] = 10'b1010011011;
    16'b0000000000001100: out_v[208] = 10'b1011001001;
    16'b0001010000010000: out_v[208] = 10'b0110101011;
    16'b0000010010001000: out_v[208] = 10'b0110011001;
    16'b0000000010011000: out_v[208] = 10'b1110010111;
    16'b0000010000001000: out_v[208] = 10'b0100010011;
    16'b0001000010010000: out_v[208] = 10'b1110010011;
    16'b0001010010011100: out_v[208] = 10'b0111001000;
    16'b0000000000001110: out_v[208] = 10'b0110010001;
    16'b0000010010011000: out_v[208] = 10'b1111111110;
    16'b0001000000011010: out_v[208] = 10'b0011110111;
    16'b0001000000010000: out_v[208] = 10'b0110110010;
    16'b0000000100001110: out_v[208] = 10'b0011111000;
    16'b0000000100001010: out_v[208] = 10'b1101101001;
    16'b0000000000000010: out_v[208] = 10'b1010100101;
    16'b0000000100000000: out_v[208] = 10'b1011110001;
    16'b0000000100000100: out_v[208] = 10'b0010001111;
    16'b0000000100000010: out_v[208] = 10'b1101000101;
    16'b0000000100000110: out_v[208] = 10'b0010011111;
    16'b0000000100001000: out_v[208] = 10'b1110111101;
    16'b0000000000001010: out_v[208] = 10'b1100100010;
    16'b0000000000000000: out_v[208] = 10'b0100100010;
    16'b0000000100001100: out_v[208] = 10'b1010011101;
    16'b0000000100011110: out_v[208] = 10'b0010001010;
    16'b0000000000000011: out_v[208] = 10'b0110101011;
    16'b0000000100010110: out_v[208] = 10'b0011010100;
    16'b0000000000000001: out_v[208] = 10'b0011001110;
    16'b0000000000010000: out_v[208] = 10'b1001010111;
    16'b0000010100000110: out_v[208] = 10'b1111001111;
    16'b0001000000001010: out_v[208] = 10'b0010011111;
    16'b0000000100000111: out_v[208] = 10'b0101000101;
    16'b0000000100000011: out_v[208] = 10'b1110111011;
    16'b0000010000000010: out_v[208] = 10'b0111000101;
    16'b0000010000010010: out_v[208] = 10'b0001010011;
    16'b0001000000000010: out_v[208] = 10'b0010111001;
    16'b0000010100010110: out_v[208] = 10'b0011101011;
    16'b0000000010000000: out_v[208] = 10'b0101010111;
    16'b0000000100001111: out_v[208] = 10'b1100111001;
    16'b0000000000001001: out_v[208] = 10'b0110100101;
    16'b0000000000001011: out_v[208] = 10'b1011100010;
    16'b0000000000011110: out_v[208] = 10'b1110011100;
    16'b0001000000011110: out_v[208] = 10'b1001100101;
    16'b0001000000001110: out_v[208] = 10'b1001000111;
    16'b0001000100001110: out_v[208] = 10'b1100010000;
    16'b0100000100001110: out_v[208] = 10'b1010111000;
    16'b0001000100011110: out_v[208] = 10'b1010110110;
    16'b0000000101001110: out_v[208] = 10'b0011101011;
    16'b0000000000000100: out_v[208] = 10'b1100011100;
    16'b0000000110001110: out_v[208] = 10'b1101110100;
    16'b0100000100011110: out_v[208] = 10'b1000111001;
    16'b0000000000000110: out_v[208] = 10'b1010111000;
    16'b0000010100011110: out_v[208] = 10'b0110001111;
    16'b0001000100000010: out_v[208] = 10'b0010111111;
    16'b0001010000010010: out_v[208] = 10'b0100010011;
    16'b0001000110001110: out_v[208] = 10'b1100100000;
    16'b0001000100000110: out_v[208] = 10'b1100001111;
    16'b0001000100010110: out_v[208] = 10'b1100110111;
    16'b0001000000010010: out_v[208] = 10'b1111101001;
    16'b0001000100001010: out_v[208] = 10'b1100001110;
    16'b0000000000010010: out_v[208] = 10'b0011010001;
    16'b0001000000000000: out_v[208] = 10'b0111110000;
    16'b0001000000000110: out_v[208] = 10'b1100110101;
    16'b0001000100010010: out_v[208] = 10'b1100011011;
    16'b0001000100011010: out_v[208] = 10'b1001010011;
    16'b0000000000010110: out_v[208] = 10'b0001011000;
    16'b0001000010000000: out_v[208] = 10'b0000110111;
    16'b0001000110000110: out_v[208] = 10'b1001010011;
    16'b0001000010001010: out_v[208] = 10'b1100001000;
    16'b0001000010001000: out_v[208] = 10'b0011101100;
    16'b0000000110000100: out_v[208] = 10'b0000110100;
    16'b0000000010001100: out_v[208] = 10'b0000111001;
    16'b0001000110001100: out_v[208] = 10'b0010110110;
    16'b0000000110001100: out_v[208] = 10'b0100110001;
    16'b0001000100001100: out_v[208] = 10'b0110001101;
    16'b0001000110000100: out_v[208] = 10'b0011100111;
    16'b0000000010000110: out_v[208] = 10'b0001110010;
    16'b0000000110000110: out_v[208] = 10'b1100101010;
    16'b0000000010000100: out_v[208] = 10'b0010101001;
    16'b0001000100000100: out_v[208] = 10'b1100100100;
    16'b0000000010001000: out_v[208] = 10'b0111101010;
    16'b0000000000010111: out_v[208] = 10'b1011101111;
    16'b0001010100010010: out_v[208] = 10'b1001100111;
    16'b0000000000000111: out_v[208] = 10'b1011000100;
    16'b0000000000000101: out_v[208] = 10'b1111001011;
    16'b0000000000001111: out_v[208] = 10'b1010111110;
    16'b0000000000001101: out_v[208] = 10'b0110011011;
    16'b0001010000000010: out_v[208] = 10'b1111111010;
    16'b0000000000010100: out_v[208] = 10'b1010110011;
    16'b0001000000010001: out_v[208] = 10'b0011101111;
    16'b0000000000010101: out_v[208] = 10'b1101110010;
    16'b0001000000010110: out_v[208] = 10'b0011011001;
    16'b0000000100001101: out_v[208] = 10'b1001100101;
    16'b0001000100010111: out_v[208] = 10'b1100011111;
    16'b0000000100010111: out_v[208] = 10'b0011111111;
    16'b0001010100010110: out_v[208] = 10'b1100110000;
    16'b0000000100010010: out_v[208] = 10'b1100111001;
    16'b0000000100011111: out_v[208] = 10'b0010000100;
    16'b0001000000010011: out_v[208] = 10'b0000011111;
    16'b0000000100000101: out_v[208] = 10'b1000111011;
    16'b0000000000010011: out_v[208] = 10'b0111100101;
    16'b0001000100011111: out_v[208] = 10'b0010110111;
    16'b0001000000011011: out_v[208] = 10'b1011100011;
    16'b0001000100010011: out_v[208] = 10'b1100110010;
    16'b0001000000000100: out_v[208] = 10'b1110001100;
    16'b0001000000100010: out_v[208] = 10'b1001110111;
    16'b0001000010000010: out_v[208] = 10'b0011111001;
    16'b0001000000100000: out_v[208] = 10'b1000111011;
    16'b0000000010001010: out_v[208] = 10'b1011000101;
    16'b0000000000100010: out_v[208] = 10'b1101101101;
    16'b0000000000011010: out_v[208] = 10'b1011101000;
    16'b0000000000100000: out_v[208] = 10'b1011100010;
    16'b0000000110001010: out_v[208] = 10'b1001101111;
    16'b0001010100011110: out_v[208] = 10'b0100100010;
    16'b0001100000000010: out_v[208] = 10'b1111001001;
    16'b0000100000000010: out_v[208] = 10'b0011110111;
    default: out_v[208] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000010000000: out_v[209] = 10'b1010101001;
    16'b0000000011000000: out_v[209] = 10'b0111010110;
    16'b1000000011000001: out_v[209] = 10'b0000000011;
    16'b0000000001000001: out_v[209] = 10'b0011110001;
    16'b1000000011000000: out_v[209] = 10'b0010000111;
    16'b1000000001000001: out_v[209] = 10'b1010001111;
    16'b0000000001010000: out_v[209] = 10'b0101001000;
    16'b1000000110000000: out_v[209] = 10'b1000110111;
    16'b0000000111000000: out_v[209] = 10'b1010110011;
    16'b0000000001000000: out_v[209] = 10'b0111011101;
    16'b0000000000000000: out_v[209] = 10'b1110001111;
    16'b1000000010000000: out_v[209] = 10'b1101111010;
    16'b1001000011000001: out_v[209] = 10'b0000000001;
    16'b1000000000000001: out_v[209] = 10'b1110001001;
    16'b0000000001010001: out_v[209] = 10'b1110100111;
    16'b0000000110000000: out_v[209] = 10'b1101001110;
    16'b1001000001000001: out_v[209] = 10'b0100010001;
    16'b0010000010000000: out_v[209] = 10'b1010111011;
    16'b1000000001000000: out_v[209] = 10'b0100111000;
    16'b0000000011000001: out_v[209] = 10'b0010010111;
    16'b1000000111000000: out_v[209] = 10'b1011101010;
    16'b1000000111000001: out_v[209] = 10'b0011001110;
    16'b1000000010000001: out_v[209] = 10'b1011100110;
    16'b0000000000010000: out_v[209] = 10'b1000001101;
    16'b0000000100000000: out_v[209] = 10'b1111010110;
    16'b0000000010010000: out_v[209] = 10'b1001100110;
    16'b0010000000000000: out_v[209] = 10'b0001000001;
    16'b0010000010010000: out_v[209] = 10'b1101001110;
    16'b0000000010000001: out_v[209] = 10'b1010001100;
    16'b0010000000010000: out_v[209] = 10'b1010110101;
    16'b1010000010010000: out_v[209] = 10'b0000110111;
    16'b1000000000000000: out_v[209] = 10'b0000101100;
    16'b1000000010010000: out_v[209] = 10'b0000111110;
    16'b1010000010000000: out_v[209] = 10'b0100011000;
    16'b1010000110000000: out_v[209] = 10'b0110110111;
    16'b1000000100000000: out_v[209] = 10'b1100101111;
    16'b1010000000000000: out_v[209] = 10'b1101001001;
    16'b0000000011010000: out_v[209] = 10'b1010110101;
    16'b1000000000010000: out_v[209] = 10'b1000011010;
    16'b0000000000000001: out_v[209] = 10'b0101100010;
    16'b0001000010000001: out_v[209] = 10'b0110010011;
    16'b0001000011000001: out_v[209] = 10'b1100111010;
    16'b0000000110000001: out_v[209] = 10'b0010110110;
    16'b0101000010000001: out_v[209] = 10'b0011110011;
    16'b0000010000000000: out_v[209] = 10'b0100101010;
    16'b0000000000100000: out_v[209] = 10'b0111100011;
    16'b0000000010100000: out_v[209] = 10'b1010100100;
    16'b0000001110000000: out_v[209] = 10'b1111101011;
    16'b0010000001000000: out_v[209] = 10'b1011000101;
    16'b0010000011000000: out_v[209] = 10'b1111001010;
    16'b0000000011010001: out_v[209] = 10'b1001010110;
    16'b0010000001010000: out_v[209] = 10'b1001010011;
    16'b0000001010000000: out_v[209] = 10'b1000101011;
    16'b0010000011010000: out_v[209] = 10'b0111000000;
    16'b0100000010000001: out_v[209] = 10'b0110010110;
    default: out_v[209] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001011000100010: out_v[210] = 10'b0100110010;
    16'b0001010010110010: out_v[210] = 10'b0011100110;
    16'b0001001010110010: out_v[210] = 10'b1111110011;
    16'b0000000000000010: out_v[210] = 10'b1001110000;
    16'b0000001000100010: out_v[210] = 10'b1100101001;
    16'b0000000010110011: out_v[210] = 10'b1000101001;
    16'b0001010010100010: out_v[210] = 10'b0110010111;
    16'b0000001010100010: out_v[210] = 10'b0001001110;
    16'b0001000010010001: out_v[210] = 10'b0110101000;
    16'b0001010000100010: out_v[210] = 10'b0001001111;
    16'b0001001000100010: out_v[210] = 10'b0011011011;
    16'b0001000000100010: out_v[210] = 10'b0100110110;
    16'b0001000000000000: out_v[210] = 10'b0110111011;
    16'b0000000010010000: out_v[210] = 10'b0011011001;
    16'b0011000010010000: out_v[210] = 10'b0100110000;
    16'b0000001001100010: out_v[210] = 10'b1011101010;
    16'b0001000010110010: out_v[210] = 10'b0000001000;
    16'b0000001010110011: out_v[210] = 10'b0111010101;
    16'b0001000010100010: out_v[210] = 10'b1010011111;
    16'b0001000010110000: out_v[210] = 10'b0001011010;
    16'b0000000010010001: out_v[210] = 10'b0110011011;
    16'b0000001011100010: out_v[210] = 10'b0101001000;
    16'b0001011001100010: out_v[210] = 10'b1100101001;
    16'b0001001001100010: out_v[210] = 10'b0010101101;
    16'b0000000000010000: out_v[210] = 10'b1110101010;
    16'b0010000000010000: out_v[210] = 10'b0001101010;
    16'b0000001011110011: out_v[210] = 10'b0011011111;
    16'b0001011010100010: out_v[210] = 10'b1000011011;
    16'b0011000010010001: out_v[210] = 10'b1111001111;
    16'b0000000000000000: out_v[210] = 10'b1101110111;
    16'b0000011011100010: out_v[210] = 10'b1110100011;
    16'b0001000000000010: out_v[210] = 10'b0101000011;
    16'b0001001010100010: out_v[210] = 10'b0001110110;
    16'b0000011001100010: out_v[210] = 10'b1001111100;
    16'b0000001010110010: out_v[210] = 10'b1100101011;
    16'b0011000000000010: out_v[210] = 10'b1011110101;
    16'b0001000010110011: out_v[210] = 10'b1110111110;
    16'b0011000000010000: out_v[210] = 10'b0100100001;
    16'b0001000010010000: out_v[210] = 10'b0000011011;
    16'b0000000010110001: out_v[210] = 10'b0100101111;
    16'b0001010010010000: out_v[210] = 10'b1110100111;
    16'b0000000010110010: out_v[210] = 10'b1101001011;
    16'b0000001011110010: out_v[210] = 10'b0101001100;
    16'b0010000010010000: out_v[210] = 10'b1001001111;
    16'b0001000010010010: out_v[210] = 10'b0101011011;
    16'b0000000010110000: out_v[210] = 10'b1111001000;
    16'b0000000000100010: out_v[210] = 10'b1100101000;
    16'b0001011011100010: out_v[210] = 10'b1010101111;
    16'b0001010001000000: out_v[210] = 10'b0000011110;
    16'b0001000001000000: out_v[210] = 10'b1011000010;
    16'b0010000001100000: out_v[210] = 10'b1101011110;
    16'b0000001001100000: out_v[210] = 10'b0110110101;
    16'b0000000001000000: out_v[210] = 10'b1010011111;
    16'b0000000001100000: out_v[210] = 10'b0111011111;
    16'b0010001001100010: out_v[210] = 10'b0010011011;
    16'b0010001001100000: out_v[210] = 10'b0011111000;
    16'b0000001000000010: out_v[210] = 10'b1111010101;
    16'b0001000001100000: out_v[210] = 10'b0110000101;
    16'b0000010001000000: out_v[210] = 10'b0001101111;
    16'b0001010000000000: out_v[210] = 10'b1100001111;
    16'b0000010000000000: out_v[210] = 10'b1011010011;
    16'b0010001000100010: out_v[210] = 10'b1011010101;
    16'b0000001001110010: out_v[210] = 10'b0110010010;
    16'b0001000001110000: out_v[210] = 10'b1001000011;
    16'b0001001001110010: out_v[210] = 10'b0011110100;
    16'b0000000001010010: out_v[210] = 10'b1010011100;
    16'b0000001000110010: out_v[210] = 10'b1100110111;
    16'b0000000011000000: out_v[210] = 10'b0000100100;
    16'b0000000001110000: out_v[210] = 10'b1111010111;
    16'b0000000001110010: out_v[210] = 10'b1100110011;
    16'b0001011001110010: out_v[210] = 10'b1011110110;
    16'b0000011001010010: out_v[210] = 10'b1110111010;
    16'b0000001001010010: out_v[210] = 10'b1011010111;
    16'b0000000011000001: out_v[210] = 10'b1100001101;
    16'b0001000001110010: out_v[210] = 10'b1000110101;
    16'b0000011001110010: out_v[210] = 10'b0111010110;
    16'b0000000001000010: out_v[210] = 10'b1100011000;
    16'b0000000001010000: out_v[210] = 10'b1100101100;
    16'b0000010001000010: out_v[210] = 10'b0001011110;
    16'b0000001001110110: out_v[210] = 10'b0010010110;
    16'b0000001011100011: out_v[210] = 10'b1100010111;
    16'b0000000000110000: out_v[210] = 10'b1100111001;
    16'b0000000000110010: out_v[210] = 10'b1100101100;
    16'b0001001011100010: out_v[210] = 10'b1001000101;
    16'b0000001001000010: out_v[210] = 10'b0110110101;
    16'b0000010001010000: out_v[210] = 10'b0010011110;
    16'b0001001000110010: out_v[210] = 10'b0101010111;
    16'b0001000001010000: out_v[210] = 10'b1101100111;
    16'b0000010001010010: out_v[210] = 10'b0011011011;
    16'b0011000000000000: out_v[210] = 10'b0000001101;
    16'b0001000000110010: out_v[210] = 10'b1101011111;
    16'b0001000000110000: out_v[210] = 10'b1011011001;
    16'b0010000000000000: out_v[210] = 10'b0100100101;
    16'b0010000000000010: out_v[210] = 10'b0010011000;
    16'b0011000000010100: out_v[210] = 10'b1010111111;
    16'b0001000000010000: out_v[210] = 10'b1001101010;
    16'b0001000010010100: out_v[210] = 10'b0111001101;
    16'b0001000000010010: out_v[210] = 10'b0101010110;
    16'b0011000000010010: out_v[210] = 10'b1011110001;
    16'b0000000011100000: out_v[210] = 10'b0110111010;
    16'b0000011000100010: out_v[210] = 10'b0001000100;
    16'b0010011000100010: out_v[210] = 10'b1011000110;
    16'b0000010001100000: out_v[210] = 10'b0100110101;
    16'b0001010001100000: out_v[210] = 10'b0111000100;
    16'b0010011001100010: out_v[210] = 10'b1111011110;
    16'b0000000000010010: out_v[210] = 10'b0110100111;
    16'b0010001000000010: out_v[210] = 10'b0110000110;
    16'b0010001001000010: out_v[210] = 10'b1101101000;
    16'b0010000001000010: out_v[210] = 10'b1101100000;
    16'b0010010000000010: out_v[210] = 10'b1001000111;
    16'b0000001000100000: out_v[210] = 10'b1110000000;
    16'b0000011001100000: out_v[210] = 10'b0001110011;
    16'b0010001000100000: out_v[210] = 10'b0101010101;
    16'b0011010000010000: out_v[210] = 10'b1010110011;
    16'b0000010000100010: out_v[210] = 10'b1011010010;
    16'b0011010010010000: out_v[210] = 10'b0010111000;
    16'b0001010000000010: out_v[210] = 10'b1100100111;
    16'b0011010000000010: out_v[210] = 10'b1111110010;
    16'b0011011001100010: out_v[210] = 10'b1000000111;
    16'b0010010000010000: out_v[210] = 10'b0111001111;
    16'b0011011000100010: out_v[210] = 10'b1111101010;
    16'b0001010000010000: out_v[210] = 10'b0111110000;
    16'b0011010000000000: out_v[210] = 10'b0001100110;
    16'b0000000001100010: out_v[210] = 10'b0111000000;
    16'b0000000000100000: out_v[210] = 10'b1010110101;
    16'b0000000011100010: out_v[210] = 10'b0011001110;
    16'b0000000011110000: out_v[210] = 10'b0111000110;
    16'b0000000011110010: out_v[210] = 10'b0010111111;
    16'b0000000010100010: out_v[210] = 10'b1001001110;
    16'b0010001011100010: out_v[210] = 10'b0010101001;
    16'b0001001001100000: out_v[210] = 10'b0001111111;
    16'b0010001100100010: out_v[210] = 10'b0110001110;
    16'b0011001000000010: out_v[210] = 10'b1110000011;
    16'b0011000001000010: out_v[210] = 10'b1110010010;
    16'b0001000001000010: out_v[210] = 10'b0010101011;
    16'b0011001001100010: out_v[210] = 10'b1001101000;
    16'b0010000001010000: out_v[210] = 10'b1110001011;
    16'b0011001001000010: out_v[210] = 10'b0111101010;
    16'b0001011001100000: out_v[210] = 10'b1101101111;
    16'b0010000001100010: out_v[210] = 10'b0111000001;
    16'b0010000001110000: out_v[210] = 10'b0110000111;
    16'b0010000001000000: out_v[210] = 10'b1000010110;
    16'b0001001001000010: out_v[210] = 10'b1111111000;
    16'b0011011001000010: out_v[210] = 10'b1110001101;
    16'b0011000001010000: out_v[210] = 10'b0111100011;
    16'b0000000100010000: out_v[210] = 10'b1001110111;
    default: out_v[210] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000001000010100: out_v[211] = 10'b0010100111;
    16'b0001001010010100: out_v[211] = 10'b0000011000;
    16'b1101001010010100: out_v[211] = 10'b0001110110;
    16'b1101011010010100: out_v[211] = 10'b0011100110;
    16'b0000001010010100: out_v[211] = 10'b1000100001;
    16'b0001001000010000: out_v[211] = 10'b0010111100;
    16'b1101001000001100: out_v[211] = 10'b0101100110;
    16'b0001011010010000: out_v[211] = 10'b0011100001;
    16'b1101001010011100: out_v[211] = 10'b0010101111;
    16'b0101001010010100: out_v[211] = 10'b1011011000;
    16'b0001001000010100: out_v[211] = 10'b0011111000;
    16'b1100001000010100: out_v[211] = 10'b1110110011;
    16'b0001011000010000: out_v[211] = 10'b1011011011;
    16'b0100001010010100: out_v[211] = 10'b1011001000;
    16'b0001001010010000: out_v[211] = 10'b0010011001;
    16'b1101000000000100: out_v[211] = 10'b0111011011;
    16'b0101001000010100: out_v[211] = 10'b0010001111;
    16'b1101001010000100: out_v[211] = 10'b0110101110;
    16'b1101000010001100: out_v[211] = 10'b1110001111;
    16'b1101001000010100: out_v[211] = 10'b0111100100;
    16'b1101000000001100: out_v[211] = 10'b0011001011;
    16'b1101001010001100: out_v[211] = 10'b0000111111;
    16'b0101001000011100: out_v[211] = 10'b1111001101;
    16'b0000000010010000: out_v[211] = 10'b1110010001;
    16'b0000001010010000: out_v[211] = 10'b1010010001;
    16'b0001011010010100: out_v[211] = 10'b0010110111;
    16'b1101001000011100: out_v[211] = 10'b1000100100;
    16'b0101011010010100: out_v[211] = 10'b1101010111;
    16'b0000000000010000: out_v[211] = 10'b0111100110;
    16'b0000001000010000: out_v[211] = 10'b0010100011;
    16'b1001001010010100: out_v[211] = 10'b0011111011;
    16'b1101000010000100: out_v[211] = 10'b0011000111;
    16'b0101001010011100: out_v[211] = 10'b1101001101;
    16'b0100001000010100: out_v[211] = 10'b0101001011;
    16'b0000000110010000: out_v[211] = 10'b0011001111;
    16'b1101011010000100: out_v[211] = 10'b0110111111;
    16'b1101001000000100: out_v[211] = 10'b0111010111;
    16'b0000000000010100: out_v[211] = 10'b0111010110;
    16'b0000001100010100: out_v[211] = 10'b1001100000;
    16'b0000000110000000: out_v[211] = 10'b0101010011;
    16'b0000000100000000: out_v[211] = 10'b1111000011;
    16'b0000000000000000: out_v[211] = 10'b1101110000;
    16'b0000000100000100: out_v[211] = 10'b0010110111;
    16'b0000000000000100: out_v[211] = 10'b0001001110;
    16'b0000000101000100: out_v[211] = 10'b1110010101;
    16'b0100000100001100: out_v[211] = 10'b1100000101;
    16'b0100000000000100: out_v[211] = 10'b0000110010;
    16'b0100000100000000: out_v[211] = 10'b1000010110;
    16'b1100000100000100: out_v[211] = 10'b0000011101;
    16'b0100000100001000: out_v[211] = 10'b0110010101;
    16'b1100000100001100: out_v[211] = 10'b0001011101;
    16'b1000000100000000: out_v[211] = 10'b0010100111;
    16'b0000000110000100: out_v[211] = 10'b1011110101;
    16'b0001000100010000: out_v[211] = 10'b0101001110;
    16'b0100010110000000: out_v[211] = 10'b1111110111;
    16'b1100000110001100: out_v[211] = 10'b1000101101;
    16'b1100000100000000: out_v[211] = 10'b1100010000;
    16'b0100000000000000: out_v[211] = 10'b0100100110;
    16'b0100000110000100: out_v[211] = 10'b1111111111;
    16'b0100000110000000: out_v[211] = 10'b0000110111;
    16'b1000000000000100: out_v[211] = 10'b0111011010;
    16'b1000000100000100: out_v[211] = 10'b0001111111;
    16'b1100000100001000: out_v[211] = 10'b0111111001;
    16'b0000000100010100: out_v[211] = 10'b0010110100;
    16'b0100000100000100: out_v[211] = 10'b1111010100;
    16'b0000000100010000: out_v[211] = 10'b0011011011;
    16'b0000010110000100: out_v[211] = 10'b0101010100;
    16'b0100010110001000: out_v[211] = 10'b1101000111;
    16'b0000010110000000: out_v[211] = 10'b0111001100;
    16'b0000010100000000: out_v[211] = 10'b1101101100;
    16'b0100000110001100: out_v[211] = 10'b0001101111;
    16'b1000000110000100: out_v[211] = 10'b1011011101;
    16'b0100010110000100: out_v[211] = 10'b1011110111;
    16'b0101000100011000: out_v[211] = 10'b1110001111;
    16'b0100000100011000: out_v[211] = 10'b1000101100;
    16'b0100000100011100: out_v[211] = 10'b1001011011;
    16'b0100000110001000: out_v[211] = 10'b1101110011;
    16'b1100000000010100: out_v[211] = 10'b1000011011;
    16'b0100010000000100: out_v[211] = 10'b0110100001;
    16'b0100010010000100: out_v[211] = 10'b1101101010;
    16'b0100000100010100: out_v[211] = 10'b0001101000;
    16'b1100000000000100: out_v[211] = 10'b0011001110;
    16'b0100000000010100: out_v[211] = 10'b1110110001;
    16'b0100001000011100: out_v[211] = 10'b1000011011;
    16'b0100001000000100: out_v[211] = 10'b0000101100;
    16'b0000000010010100: out_v[211] = 10'b1111100011;
    16'b0000000010000100: out_v[211] = 10'b0010100010;
    16'b1100000000001100: out_v[211] = 10'b0000100111;
    16'b0000001000000100: out_v[211] = 10'b1010001110;
    16'b1000000100010100: out_v[211] = 10'b0011001101;
    16'b0000010010000100: out_v[211] = 10'b1011011111;
    16'b0000010010000000: out_v[211] = 10'b0011001010;
    16'b0000000110010100: out_v[211] = 10'b0010111011;
    16'b0100000000001100: out_v[211] = 10'b1110111010;
    16'b0000000010000000: out_v[211] = 10'b0000111110;
    16'b0100001000001100: out_v[211] = 10'b1111011010;
    16'b1100000100010100: out_v[211] = 10'b0010011101;
    16'b1100000110000100: out_v[211] = 10'b1001011011;
    16'b0100000010000100: out_v[211] = 10'b1001101011;
    16'b1001001100010100: out_v[211] = 10'b1001011011;
    16'b0001001110010000: out_v[211] = 10'b1011000100;
    16'b1001001000010100: out_v[211] = 10'b0010011100;
    16'b0001001100010000: out_v[211] = 10'b0001111000;
    16'b0000001110010000: out_v[211] = 10'b1100000011;
    16'b1001001110010100: out_v[211] = 10'b1000110011;
    16'b1000001000010000: out_v[211] = 10'b0000110111;
    16'b1001001100010000: out_v[211] = 10'b1000111111;
    16'b0001001100010100: out_v[211] = 10'b0011011111;
    16'b0000001100010000: out_v[211] = 10'b1001010000;
    16'b1101001110010100: out_v[211] = 10'b1011000011;
    16'b1001000100010100: out_v[211] = 10'b1101100010;
    16'b1000001100010100: out_v[211] = 10'b0100110111;
    16'b0001001110010100: out_v[211] = 10'b1100101111;
    16'b1101001100010100: out_v[211] = 10'b1100010011;
    16'b1000001000010100: out_v[211] = 10'b1011000001;
    16'b1001001110010000: out_v[211] = 10'b0011010101;
    16'b1001000100000100: out_v[211] = 10'b1000110011;
    16'b1001001000010000: out_v[211] = 10'b1001001000;
    16'b1000001100010000: out_v[211] = 10'b1101101000;
    16'b1100001010010100: out_v[211] = 10'b1110010111;
    16'b1000001010010100: out_v[211] = 10'b1101100110;
    16'b0100001100010100: out_v[211] = 10'b1011100101;
    16'b0000001010000000: out_v[211] = 10'b1000111000;
    16'b0000001110010100: out_v[211] = 10'b0110100100;
    16'b0000001000000000: out_v[211] = 10'b0010011011;
    16'b1100001100010100: out_v[211] = 10'b0011110001;
    16'b1000001000000100: out_v[211] = 10'b0000111110;
    16'b1100001000000100: out_v[211] = 10'b1111110111;
    16'b1100001010000100: out_v[211] = 10'b1110100001;
    16'b1000001110010100: out_v[211] = 10'b0110000010;
    16'b1000001010000100: out_v[211] = 10'b1001100110;
    16'b0000001010000100: out_v[211] = 10'b0011011110;
    16'b1100001000001100: out_v[211] = 10'b0000111000;
    16'b1101001100011100: out_v[211] = 10'b1101101010;
    16'b0101001100010000: out_v[211] = 10'b0111010110;
    16'b0101001100010100: out_v[211] = 10'b1111001110;
    16'b1101001100010000: out_v[211] = 10'b1001001000;
    16'b0101001100011100: out_v[211] = 10'b1000111011;
    16'b0100001100010000: out_v[211] = 10'b1001111011;
    16'b0101001000010000: out_v[211] = 10'b1011011011;
    16'b1100001100011100: out_v[211] = 10'b1101110010;
    16'b0100001000010000: out_v[211] = 10'b1000111000;
    16'b0100001100011100: out_v[211] = 10'b0001110011;
    16'b1000001010000000: out_v[211] = 10'b1011010110;
    16'b1000000010000000: out_v[211] = 10'b1100010011;
    16'b1000000000000000: out_v[211] = 10'b0101110001;
    16'b1000000100010000: out_v[211] = 10'b0110000111;
    16'b1000001000000000: out_v[211] = 10'b1001010111;
    16'b1000000110000000: out_v[211] = 10'b0011010100;
    16'b0001001000000000: out_v[211] = 10'b0111101011;
    16'b1001001000000100: out_v[211] = 10'b1101101011;
    16'b1001001000000000: out_v[211] = 10'b0011101011;
    16'b1001001010010000: out_v[211] = 10'b1101101111;
    16'b1001000000000100: out_v[211] = 10'b1111001100;
    16'b1001001010000000: out_v[211] = 10'b0000100111;
    16'b0000001110000000: out_v[211] = 10'b0110001110;
    16'b0000001110000100: out_v[211] = 10'b0111011101;
    16'b0000001100000100: out_v[211] = 10'b0110000011;
    16'b1000001110010000: out_v[211] = 10'b0100011110;
    16'b1100001110000100: out_v[211] = 10'b1111000001;
    16'b1000001100000100: out_v[211] = 10'b0110000001;
    16'b0000001100000000: out_v[211] = 10'b0110001100;
    16'b1000001100000000: out_v[211] = 10'b0110001111;
    16'b1100001110010100: out_v[211] = 10'b1111010010;
    16'b1000001110000100: out_v[211] = 10'b1111000111;
    16'b1100001100000000: out_v[211] = 10'b0100001110;
    16'b1100001100000100: out_v[211] = 10'b0110010011;
    16'b1000001110000000: out_v[211] = 10'b0011100000;
    16'b1001001100000100: out_v[211] = 10'b1001101010;
    16'b0001001100000000: out_v[211] = 10'b1011011101;
    16'b1001000000010100: out_v[211] = 10'b1011100011;
    16'b1001000100010000: out_v[211] = 10'b1100110110;
    16'b1101000100010100: out_v[211] = 10'b1101010100;
    default: out_v[211] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100000001000000: out_v[212] = 10'b1100101110;
    16'b0100010101010000: out_v[212] = 10'b0101010101;
    16'b0110110111010010: out_v[212] = 10'b1011111001;
    16'b0100110011010010: out_v[212] = 10'b0100111101;
    16'b0000010001000010: out_v[212] = 10'b1001011011;
    16'b0100000001010010: out_v[212] = 10'b0111001010;
    16'b0110110010010000: out_v[212] = 10'b1001001000;
    16'b0100000001000010: out_v[212] = 10'b0111000001;
    16'b0100110001010000: out_v[212] = 10'b0100011110;
    16'b0110010010010010: out_v[212] = 10'b1011100011;
    16'b0100000001010000: out_v[212] = 10'b1101010010;
    16'b0100000101010000: out_v[212] = 10'b1001111011;
    16'b0100000101000000: out_v[212] = 10'b0111110110;
    16'b0000010001010000: out_v[212] = 10'b0111100110;
    16'b0100010001010000: out_v[212] = 10'b0110110001;
    16'b0100010001000000: out_v[212] = 10'b1011111100;
    16'b0100110101010000: out_v[212] = 10'b0110000010;
    16'b0100110010010010: out_v[212] = 10'b0101011011;
    16'b0100010001000010: out_v[212] = 10'b0001111001;
    16'b0100110001010010: out_v[212] = 10'b0110101011;
    16'b0110110011010010: out_v[212] = 10'b0100010111;
    16'b0110110010010010: out_v[212] = 10'b1111101011;
    16'b0100010001010010: out_v[212] = 10'b1101101010;
    16'b0010110010010010: out_v[212] = 10'b0110111111;
    16'b0100010010010010: out_v[212] = 10'b0101110111;
    16'b0100010011010010: out_v[212] = 10'b1000111001;
    16'b0110110110010000: out_v[212] = 10'b1101110011;
    16'b0000010001010010: out_v[212] = 10'b0001001111;
    16'b0000000001000010: out_v[212] = 10'b0101010010;
    16'b0100110111010000: out_v[212] = 10'b1111000011;
    16'b0100100011010010: out_v[212] = 10'b0111001000;
    16'b0000010001000000: out_v[212] = 10'b1000111001;
    16'b0100110111010010: out_v[212] = 10'b1011110101;
    16'b0100110110010000: out_v[212] = 10'b0001010111;
    16'b0000110010010010: out_v[212] = 10'b1101001011;
    16'b0100010101000000: out_v[212] = 10'b1000111110;
    16'b0000010011010010: out_v[212] = 10'b0011001110;
    16'b0100110010010000: out_v[212] = 10'b1110000111;
    16'b0100010111010000: out_v[212] = 10'b0110111110;
    16'b0100000000000010: out_v[212] = 10'b0010010111;
    16'b0110010011010010: out_v[212] = 10'b1110101011;
    16'b0000000001000000: out_v[212] = 10'b0000010001;
    16'b0100010101010010: out_v[212] = 10'b0100111010;
    16'b0000110010010000: out_v[212] = 10'b1111111010;
    16'b0000010010010000: out_v[212] = 10'b0111001110;
    16'b0100110011010000: out_v[212] = 10'b1000100110;
    16'b0100010011010000: out_v[212] = 10'b1011111110;
    16'b0000000000000010: out_v[212] = 10'b1110000101;
    16'b0000000100000010: out_v[212] = 10'b0011010111;
    16'b0100000000000000: out_v[212] = 10'b1110011001;
    16'b0000000000000000: out_v[212] = 10'b0111100010;
    16'b0000000000010010: out_v[212] = 10'b1010101011;
    16'b0100000100000010: out_v[212] = 10'b1011100010;
    16'b0000000000010000: out_v[212] = 10'b1010100100;
    16'b0000010000010010: out_v[212] = 10'b1000110110;
    16'b0000010000010000: out_v[212] = 10'b0000110111;
    16'b0100000000010010: out_v[212] = 10'b0010110110;
    16'b0100000000000110: out_v[212] = 10'b0000011110;
    16'b0000000001010110: out_v[212] = 10'b1000110101;
    16'b0000000000000110: out_v[212] = 10'b1100110100;
    16'b0000000000010110: out_v[212] = 10'b1111100000;
    16'b0000110011010010: out_v[212] = 10'b0111010101;
    16'b0000110000010010: out_v[212] = 10'b1001011010;
    16'b0000000001010010: out_v[212] = 10'b1101100110;
    16'b0100110000010010: out_v[212] = 10'b0000011110;
    16'b0100010000010010: out_v[212] = 10'b0100011100;
    16'b0000110000010110: out_v[212] = 10'b0000111110;
    16'b0000100001010110: out_v[212] = 10'b1010101110;
    16'b0100000000010110: out_v[212] = 10'b1110011010;
    16'b0000100000010010: out_v[212] = 10'b1101101100;
    16'b0000100000010110: out_v[212] = 10'b1111110101;
    16'b0000100000010000: out_v[212] = 10'b0010111101;
    16'b0100100000010010: out_v[212] = 10'b1010110000;
    16'b0100110000010000: out_v[212] = 10'b0101011010;
    16'b0100100000010000: out_v[212] = 10'b0001100111;
    16'b0000100001010010: out_v[212] = 10'b0101110110;
    16'b0000110001010010: out_v[212] = 10'b1111011000;
    16'b0100100001010010: out_v[212] = 10'b0011100001;
    16'b0000110000010000: out_v[212] = 10'b1000101111;
    16'b0100000000010000: out_v[212] = 10'b1100011110;
    16'b0110000000000010: out_v[212] = 10'b1000000110;
    16'b0110000000010010: out_v[212] = 10'b0000010111;
    16'b0000000101000000: out_v[212] = 10'b1011011100;
    16'b0100000100000000: out_v[212] = 10'b0101011011;
    16'b0100010100000000: out_v[212] = 10'b1100111110;
    16'b0000000100000000: out_v[212] = 10'b0000100110;
    16'b0000100001010000: out_v[212] = 10'b0100110110;
    16'b0000000101010000: out_v[212] = 10'b0101110001;
    16'b0000000001010000: out_v[212] = 10'b0010100101;
    16'b0000000100010000: out_v[212] = 10'b1011110111;
    16'b0100000100010000: out_v[212] = 10'b1101100000;
    16'b0000010101000000: out_v[212] = 10'b0111001101;
    16'b0100000101000010: out_v[212] = 10'b1010000100;
    16'b0100110100010000: out_v[212] = 10'b0011010110;
    16'b0100010100010000: out_v[212] = 10'b1000010101;
    16'b0100000000001000: out_v[212] = 10'b0111111000;
    16'b0000010010000000: out_v[212] = 10'b0010110000;
    16'b0000000011000000: out_v[212] = 10'b0000111111;
    16'b0000000011000010: out_v[212] = 10'b1011010010;
    16'b0100010111000010: out_v[212] = 10'b1111110010;
    16'b0000000010000000: out_v[212] = 10'b1011010000;
    16'b0000000101000010: out_v[212] = 10'b0101011000;
    16'b0100010101000010: out_v[212] = 10'b1010010011;
    16'b0000010101000010: out_v[212] = 10'b1110101010;
    16'b0000010111000010: out_v[212] = 10'b0011011110;
    16'b0100000011000000: out_v[212] = 10'b1010110100;
    16'b0000010011000010: out_v[212] = 10'b1100110011;
    16'b0000010011000000: out_v[212] = 10'b0100011011;
    16'b0000000001001000: out_v[212] = 10'b0001110111;
    16'b0000001001001000: out_v[212] = 10'b1011111011;
    16'b0100010011000000: out_v[212] = 10'b1001111011;
    16'b0000001011001000: out_v[212] = 10'b0010101101;
    16'b0000000011001000: out_v[212] = 10'b0000011111;
    16'b0100010011000010: out_v[212] = 10'b0000111001;
    16'b0100000111000000: out_v[212] = 10'b0001111101;
    16'b0100100001010000: out_v[212] = 10'b0010111100;
    16'b0000000001000110: out_v[212] = 10'b1011000001;
    16'b0010000011000010: out_v[212] = 10'b1010011011;
    16'b0010000001000010: out_v[212] = 10'b1001110010;
    16'b0100000001000110: out_v[212] = 10'b1110110111;
    16'b0010000010000010: out_v[212] = 10'b1011001000;
    16'b0010000001000110: out_v[212] = 10'b1110111111;
    16'b0010000011000110: out_v[212] = 10'b1110111100;
    16'b0100000011010010: out_v[212] = 10'b0110001110;
    16'b0100000011000010: out_v[212] = 10'b0110111111;
    16'b0100010100000010: out_v[212] = 10'b0100011000;
    16'b0100010000000000: out_v[212] = 10'b1100101101;
    16'b0100001000001000: out_v[212] = 10'b0110110001;
    16'b0100010110000010: out_v[212] = 10'b1001111010;
    16'b0100010100100010: out_v[212] = 10'b1101101111;
    16'b0100000001001000: out_v[212] = 10'b1001001111;
    16'b0100010000001000: out_v[212] = 10'b1111110011;
    16'b0100010000000010: out_v[212] = 10'b1001110111;
    16'b0000010000000000: out_v[212] = 10'b1010100011;
    16'b0000010100000010: out_v[212] = 10'b1110000111;
    16'b0100010000100010: out_v[212] = 10'b0011110011;
    16'b0100010010000000: out_v[212] = 10'b1101000010;
    16'b0100000010000000: out_v[212] = 10'b1111101010;
    16'b0100010100010010: out_v[212] = 10'b1111000100;
    16'b0000010000000010: out_v[212] = 10'b0111101001;
    16'b0100010000010000: out_v[212] = 10'b0011110001;
    16'b0000010100010000: out_v[212] = 10'b0101010101;
    16'b0000010100000000: out_v[212] = 10'b0001000110;
    16'b0100000011001000: out_v[212] = 10'b1101101110;
    16'b0100001010001000: out_v[212] = 10'b1111100111;
    16'b0100001001001000: out_v[212] = 10'b1000001010;
    16'b0100001011001000: out_v[212] = 10'b0110011001;
    16'b0100000010001000: out_v[212] = 10'b1111010101;
    16'b0100010010001000: out_v[212] = 10'b1000101111;
    16'b0100010011001000: out_v[212] = 10'b0011110101;
    default: out_v[212] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000011101000: out_v[213] = 10'b0010110100;
    16'b0010011011101001: out_v[213] = 10'b1011011011;
    16'b0010000011101010: out_v[213] = 10'b0110111011;
    16'b0010001011101000: out_v[213] = 10'b1110100010;
    16'b0000011011000001: out_v[213] = 10'b0100101001;
    16'b0010000010101000: out_v[213] = 10'b1101001011;
    16'b0000011011101000: out_v[213] = 10'b0110100101;
    16'b0000011011001001: out_v[213] = 10'b1101111010;
    16'b0010000011001001: out_v[213] = 10'b0010101010;
    16'b0000011001001001: out_v[213] = 10'b1000101111;
    16'b0010000011101001: out_v[213] = 10'b1011110100;
    16'b0010000011100000: out_v[213] = 10'b1011001111;
    16'b0010011011101011: out_v[213] = 10'b0001010001;
    16'b0000011011101001: out_v[213] = 10'b1001101110;
    16'b0000011011011001: out_v[213] = 10'b1001000101;
    16'b0010000011101000: out_v[213] = 10'b0000110001;
    16'b0010001011001001: out_v[213] = 10'b1100011000;
    16'b0000010011101000: out_v[213] = 10'b1000011111;
    16'b0000001011001001: out_v[213] = 10'b1011101011;
    16'b0000011011101011: out_v[213] = 10'b1110011011;
    16'b0001011011101000: out_v[213] = 10'b1010011101;
    16'b0010011011011001: out_v[213] = 10'b1010110011;
    16'b0010000011001000: out_v[213] = 10'b0100110101;
    16'b0010011011101000: out_v[213] = 10'b0111111110;
    16'b0010001011101011: out_v[213] = 10'b1001010001;
    16'b0000011011001011: out_v[213] = 10'b0100110010;
    16'b0000011010001001: out_v[213] = 10'b1100010001;
    16'b0010000011001011: out_v[213] = 10'b0011111111;
    16'b0010001011101001: out_v[213] = 10'b1011001111;
    16'b0010000001101010: out_v[213] = 10'b0001001101;
    16'b0010011011001001: out_v[213] = 10'b1111101001;
    16'b0000010011001001: out_v[213] = 10'b1011010111;
    16'b0000000011001001: out_v[213] = 10'b1011100111;
    16'b0000011010101000: out_v[213] = 10'b0101111111;
    16'b0000000010001010: out_v[213] = 10'b1010001000;
    16'b0000000000100000: out_v[213] = 10'b0010110111;
    16'b0000000000000000: out_v[213] = 10'b0001101011;
    16'b0000000000101000: out_v[213] = 10'b1111011101;
    16'b0000000000001000: out_v[213] = 10'b0110010011;
    16'b0000000010001000: out_v[213] = 10'b0010100110;
    16'b0000000010000010: out_v[213] = 10'b0010011111;
    16'b0000000011000010: out_v[213] = 10'b0001001011;
    16'b0000000000110001: out_v[213] = 10'b1001000111;
    16'b0000000000101010: out_v[213] = 10'b0000100011;
    16'b0000000000001010: out_v[213] = 10'b1101100011;
    16'b0000000011001010: out_v[213] = 10'b0010011010;
    16'b0000000010101010: out_v[213] = 10'b0111001100;
    16'b0000000000100001: out_v[213] = 10'b1011110010;
    16'b0000000000101001: out_v[213] = 10'b1001010011;
    16'b0000000000011011: out_v[213] = 10'b0011111010;
    16'b0000000001101011: out_v[213] = 10'b1010011001;
    16'b0010010011101000: out_v[213] = 10'b1001100110;
    16'b0000000000101011: out_v[213] = 10'b0000101110;
    16'b0000000000001011: out_v[213] = 10'b0101001101;
    16'b0010000011000000: out_v[213] = 10'b0110000111;
    16'b0000000011101011: out_v[213] = 10'b1011001101;
    16'b0010000001101000: out_v[213] = 10'b0110111111;
    16'b0000000000111011: out_v[213] = 10'b1011001100;
    16'b0000000011100010: out_v[213] = 10'b1111011101;
    16'b0000000011010011: out_v[213] = 10'b1101000110;
    16'b0000000001001010: out_v[213] = 10'b1101001101;
    16'b0000000001111011: out_v[213] = 10'b0011110101;
    16'b0000000011000011: out_v[213] = 10'b1110001100;
    16'b0010000011100011: out_v[213] = 10'b0100011110;
    16'b0000000001101010: out_v[213] = 10'b0010110101;
    16'b0010010011100000: out_v[213] = 10'b1001011110;
    16'b0010000011100001: out_v[213] = 10'b0110011110;
    16'b0010000011111001: out_v[213] = 10'b0011100010;
    16'b0010000011100010: out_v[213] = 10'b1000001110;
    16'b0000010001001010: out_v[213] = 10'b1001001111;
    16'b0010000001101011: out_v[213] = 10'b1010010100;
    16'b0010000011101011: out_v[213] = 10'b1110100110;
    16'b0000000011101010: out_v[213] = 10'b0111011000;
    16'b0000000011001011: out_v[213] = 10'b0110000011;
    16'b0000000011111011: out_v[213] = 10'b1011110111;
    16'b0000000001101001: out_v[213] = 10'b0000110011;
    16'b0010010011101010: out_v[213] = 10'b1101011100;
    16'b0000000011100011: out_v[213] = 10'b0110001101;
    16'b0010000011001010: out_v[213] = 10'b1011110010;
    16'b0000010001101010: out_v[213] = 10'b0010110010;
    16'b0000000011011011: out_v[213] = 10'b0111000110;
    16'b0010000011111011: out_v[213] = 10'b0101110111;
    16'b0000000010000011: out_v[213] = 10'b1001001110;
    16'b0000000001001011: out_v[213] = 10'b1110100011;
    16'b0010000010100000: out_v[213] = 10'b1100000111;
    16'b0000010011101010: out_v[213] = 10'b1010101111;
    16'b0010010001101010: out_v[213] = 10'b1001110110;
    16'b0010000000001011: out_v[213] = 10'b0101110101;
    16'b0000000000001001: out_v[213] = 10'b0111001100;
    16'b0010000010000011: out_v[213] = 10'b1111010001;
    16'b0010000010101010: out_v[213] = 10'b1000100100;
    16'b0000000010100010: out_v[213] = 10'b0101011011;
    16'b0000000000011001: out_v[213] = 10'b0110110000;
    16'b0010010000011011: out_v[213] = 10'b1111001001;
    16'b0010000000101010: out_v[213] = 10'b1000000111;
    16'b0000000010001001: out_v[213] = 10'b1001100011;
    16'b0010010010001011: out_v[213] = 10'b0101111110;
    16'b0010000010101011: out_v[213] = 10'b0001011101;
    16'b0000000010101011: out_v[213] = 10'b1100000011;
    16'b0000000001001001: out_v[213] = 10'b0011001111;
    16'b0010000010001011: out_v[213] = 10'b1001110011;
    16'b0000000010011011: out_v[213] = 10'b0110010111;
    16'b0000000010001011: out_v[213] = 10'b0101010111;
    16'b0000000000010001: out_v[213] = 10'b1011010011;
    16'b0010000001001011: out_v[213] = 10'b0011001011;
    16'b0010000010100010: out_v[213] = 10'b0001110110;
    16'b0010010011001011: out_v[213] = 10'b0011100011;
    16'b0010010000001011: out_v[213] = 10'b1000001100;
    16'b0000000000000001: out_v[213] = 10'b0111001000;
    16'b0010001010000011: out_v[213] = 10'b1101010111;
    16'b0010001000100000: out_v[213] = 10'b0101011001;
    16'b0000001000011011: out_v[213] = 10'b1011100111;
    16'b0000011010000010: out_v[213] = 10'b1000111010;
    16'b0011001000100000: out_v[213] = 10'b0010011001;
    16'b0000001010100010: out_v[213] = 10'b0011101101;
    16'b0010000010000010: out_v[213] = 10'b0000011001;
    16'b0010001010100010: out_v[213] = 10'b0001011010;
    16'b0010001000100010: out_v[213] = 10'b0010111010;
    16'b0010000000100000: out_v[213] = 10'b0111011100;
    16'b0010000000100010: out_v[213] = 10'b0011100001;
    16'b0010001000000001: out_v[213] = 10'b0011111010;
    16'b0010000000000000: out_v[213] = 10'b1010000010;
    16'b0000000000100010: out_v[213] = 10'b1110110100;
    16'b0000001010000010: out_v[213] = 10'b1000111011;
    16'b0010001010010011: out_v[213] = 10'b0101010111;
    16'b0010001010010001: out_v[213] = 10'b0111011010;
    16'b0000010010100010: out_v[213] = 10'b1111101110;
    16'b0000000000000010: out_v[213] = 10'b1000011101;
    16'b0010001000011011: out_v[213] = 10'b0111010110;
    16'b0010001010100000: out_v[213] = 10'b1101111010;
    16'b0010001010011011: out_v[213] = 10'b1110001001;
    16'b0000011010100010: out_v[213] = 10'b1100111111;
    16'b0000001000101010: out_v[213] = 10'b0010110111;
    16'b0010001000010011: out_v[213] = 10'b1001100111;
    16'b0010011010100010: out_v[213] = 10'b0100110110;
    16'b0010001010100011: out_v[213] = 10'b1001101101;
    16'b0001000011101000: out_v[213] = 10'b1011111011;
    16'b0001000011100000: out_v[213] = 10'b1011001010;
    16'b0001000001100010: out_v[213] = 10'b1110001111;
    16'b0000000010101001: out_v[213] = 10'b0110111101;
    16'b0001001010101000: out_v[213] = 10'b0011011111;
    16'b0000000010101000: out_v[213] = 10'b0110100100;
    16'b0001000010100000: out_v[213] = 10'b0001111001;
    16'b0001000010101000: out_v[213] = 10'b0011110111;
    16'b0000000011101001: out_v[213] = 10'b1001110000;
    16'b0000000010011001: out_v[213] = 10'b0011100111;
    16'b0000000011100000: out_v[213] = 10'b0100111001;
    16'b0001000001000010: out_v[213] = 10'b1011110000;
    16'b0000000001000010: out_v[213] = 10'b0000110001;
    16'b0001000001100000: out_v[213] = 10'b0010100000;
    16'b0000001010001001: out_v[213] = 10'b1111001101;
    16'b0000000001100010: out_v[213] = 10'b1111110000;
    16'b0000000001000001: out_v[213] = 10'b1011101110;
    16'b0000000010100000: out_v[213] = 10'b1101100101;
    16'b0001000000100000: out_v[213] = 10'b1100100101;
    16'b0001000000100010: out_v[213] = 10'b1000101110;
    16'b0000001010011001: out_v[213] = 10'b1010000111;
    16'b0000000001100000: out_v[213] = 10'b0100001011;
    16'b0010000000000011: out_v[213] = 10'b1000100101;
    16'b0000000001101000: out_v[213] = 10'b0111011110;
    16'b0010000001100000: out_v[213] = 10'b1110011000;
    16'b0010011001100011: out_v[213] = 10'b0111110110;
    16'b0010011000100001: out_v[213] = 10'b1111101111;
    16'b0010010001100000: out_v[213] = 10'b1001001010;
    16'b0010010000100000: out_v[213] = 10'b1000101011;
    16'b0010000000100011: out_v[213] = 10'b1011000111;
    16'b0010000000101000: out_v[213] = 10'b0110011000;
    16'b0010010001100001: out_v[213] = 10'b1110101010;
    16'b0010011001100010: out_v[213] = 10'b1100101011;
    16'b0010011001100000: out_v[213] = 10'b1111000000;
    16'b0010011000100000: out_v[213] = 10'b0011101110;
    16'b0010000000000001: out_v[213] = 10'b1101101010;
    16'b0010000000100001: out_v[213] = 10'b1111010101;
    16'b0010011001100001: out_v[213] = 10'b1000011110;
    16'b0010010000000001: out_v[213] = 10'b1011110011;
    16'b0010000001100010: out_v[213] = 10'b0101100010;
    16'b0010010001101000: out_v[213] = 10'b1011010011;
    16'b0000011001100010: out_v[213] = 10'b0111101011;
    16'b0000011001100011: out_v[213] = 10'b1001111000;
    16'b0000010001100000: out_v[213] = 10'b1100001110;
    16'b0010011000100011: out_v[213] = 10'b0011101111;
    16'b0010010000100001: out_v[213] = 10'b1111001000;
    16'b0010010000100011: out_v[213] = 10'b1001111000;
    16'b0010010001100010: out_v[213] = 10'b0100000101;
    16'b0010010001100011: out_v[213] = 10'b1110110011;
    16'b0010001010101010: out_v[213] = 10'b1001101100;
    16'b0010000010001010: out_v[213] = 10'b1000100101;
    16'b0010001000101010: out_v[213] = 10'b1101101110;
    16'b0010000000000010: out_v[213] = 10'b1011100010;
    16'b0010001010101000: out_v[213] = 10'b1001000010;
    16'b0000001010101010: out_v[213] = 10'b1011001011;
    16'b0010001100000011: out_v[213] = 10'b1001111011;
    16'b0010000010001000: out_v[213] = 10'b1101000100;
    16'b0000001000100010: out_v[213] = 10'b1101100111;
    16'b0010001000000011: out_v[213] = 10'b1110000110;
    16'b0011000011101010: out_v[213] = 10'b1111110010;
    16'b0011000011101000: out_v[213] = 10'b1111000111;
    16'b0000000000000011: out_v[213] = 10'b1110100111;
    16'b0001000011101010: out_v[213] = 10'b0111010100;
    16'b0000001010011011: out_v[213] = 10'b0111011110;
    16'b0001000011001010: out_v[213] = 10'b0111010001;
    16'b0000001010001011: out_v[213] = 10'b0110010100;
    16'b0011000011001000: out_v[213] = 10'b0101001011;
    16'b0010001000101011: out_v[213] = 10'b1001000111;
    16'b0010001000101000: out_v[213] = 10'b0101010010;
    16'b0000001000001011: out_v[213] = 10'b0101111011;
    16'b0010001000001011: out_v[213] = 10'b0001110111;
    16'b0000001000010011: out_v[213] = 10'b1100100001;
    16'b0010001010101011: out_v[213] = 10'b1011101001;
    default: out_v[213] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000010011100: out_v[214] = 10'b0001000111;
    16'b0001001010001000: out_v[214] = 10'b0010011101;
    16'b0001011010001100: out_v[214] = 10'b0110000111;
    16'b0001011010011100: out_v[214] = 10'b1100110111;
    16'b0000001010001000: out_v[214] = 10'b1110010000;
    16'b0001011010001000: out_v[214] = 10'b1001101111;
    16'b0001010010011100: out_v[214] = 10'b0001001100;
    16'b0000000010011000: out_v[214] = 10'b0100110011;
    16'b0000001010001100: out_v[214] = 10'b0011110011;
    16'b0001000010011100: out_v[214] = 10'b0111110110;
    16'b0000000010001000: out_v[214] = 10'b1101001100;
    16'b0000000010010100: out_v[214] = 10'b1010100111;
    16'b0000000010001100: out_v[214] = 10'b0010000001;
    16'b0000001010011000: out_v[214] = 10'b0111000101;
    16'b0001010000011100: out_v[214] = 10'b0010111100;
    16'b0001010000010100: out_v[214] = 10'b0000100001;
    16'b0000010010011100: out_v[214] = 10'b0111011110;
    16'b0000001000000000: out_v[214] = 10'b1111100111;
    16'b0000001000011000: out_v[214] = 10'b1001111100;
    16'b0000001010011100: out_v[214] = 10'b1010100011;
    16'b0000000000000000: out_v[214] = 10'b0110110011;
    16'b0001001010011000: out_v[214] = 10'b0111011011;
    16'b0000001000001000: out_v[214] = 10'b1011001000;
    16'b0001001010000000: out_v[214] = 10'b1001010011;
    16'b0001001010011100: out_v[214] = 10'b0111101100;
    16'b0000010000010100: out_v[214] = 10'b0110101011;
    16'b0000000000011100: out_v[214] = 10'b0100100011;
    16'b0000000000010100: out_v[214] = 10'b1000001100;
    16'b0001010010001100: out_v[214] = 10'b0111010010;
    16'b0001011000011100: out_v[214] = 10'b0100000011;
    16'b0000000000011000: out_v[214] = 10'b0101110101;
    16'b0001011010011000: out_v[214] = 10'b1111111011;
    16'b0001001011001000: out_v[214] = 10'b1101111011;
    16'b0000000000001100: out_v[214] = 10'b0010100110;
    16'b0000101000000000: out_v[214] = 10'b1101110010;
    16'b0000101000010000: out_v[214] = 10'b0010001001;
    16'b0000100000000000: out_v[214] = 10'b0001010011;
    16'b0000101000011000: out_v[214] = 10'b0001011010;
    16'b0000101000011100: out_v[214] = 10'b0001010111;
    16'b0010100000000000: out_v[214] = 10'b0101010011;
    16'b0110100000000000: out_v[214] = 10'b1001100110;
    16'b0000001000010000: out_v[214] = 10'b1110001100;
    16'b0000101000010100: out_v[214] = 10'b0000111100;
    16'b0000001000011100: out_v[214] = 10'b0000111100;
    16'b0000100000010100: out_v[214] = 10'b1000001010;
    16'b0000101000000100: out_v[214] = 10'b0011110101;
    16'b0000100000010000: out_v[214] = 10'b1011000100;
    16'b0000100000001000: out_v[214] = 10'b1110001100;
    16'b0000001000010100: out_v[214] = 10'b1101011010;
    16'b0000101000001000: out_v[214] = 10'b0110000001;
    16'b0000101001010100: out_v[214] = 10'b0001101010;
    16'b0000100000011100: out_v[214] = 10'b1000111011;
    16'b0000111000010000: out_v[214] = 10'b1000100111;
    16'b0000111000011000: out_v[214] = 10'b1011100111;
    16'b0000101010011000: out_v[214] = 10'b1001110101;
    16'b0000101001011000: out_v[214] = 10'b0101000001;
    16'b0000101000001100: out_v[214] = 10'b0010001110;
    16'b0000101001010000: out_v[214] = 10'b1111010111;
    16'b0000101001000100: out_v[214] = 10'b0110000111;
    16'b0000100000000100: out_v[214] = 10'b0011111000;
    16'b0000001000000100: out_v[214] = 10'b1110110110;
    16'b0000101001011100: out_v[214] = 10'b1011011101;
    16'b0000101001000000: out_v[214] = 10'b1110001110;
    16'b0000100000011000: out_v[214] = 10'b0100111110;
    16'b0000101010011100: out_v[214] = 10'b0111100000;
    16'b0000000000010000: out_v[214] = 10'b0100001001;
    16'b0000100010011100: out_v[214] = 10'b1011000100;
    16'b0000000001010100: out_v[214] = 10'b0010101001;
    16'b0010000001010100: out_v[214] = 10'b1011011110;
    16'b0010001001010000: out_v[214] = 10'b1000110111;
    16'b0000000010000100: out_v[214] = 10'b0111011001;
    16'b0000001010010100: out_v[214] = 10'b1011101101;
    16'b0000000000000100: out_v[214] = 10'b1001111001;
    16'b0000001001000000: out_v[214] = 10'b1110111001;
    16'b0000001001010000: out_v[214] = 10'b1001111011;
    16'b0110000000010100: out_v[214] = 10'b1111010001;
    16'b0000000010010000: out_v[214] = 10'b1000001010;
    16'b0000100010010100: out_v[214] = 10'b1110100011;
    16'b0000010010010100: out_v[214] = 10'b1001101010;
    16'b0000100010001100: out_v[214] = 10'b1101001101;
    16'b0000100010000100: out_v[214] = 10'b0111111011;
    16'b0000111010001000: out_v[214] = 10'b0111110010;
    16'b0000101010000000: out_v[214] = 10'b0011100010;
    16'b0000100010011000: out_v[214] = 10'b1000110110;
    16'b0000101010001000: out_v[214] = 10'b1101001101;
    16'b0000001010000000: out_v[214] = 10'b0100110110;
    16'b0000000010000000: out_v[214] = 10'b0111110101;
    16'b0000101010000100: out_v[214] = 10'b0000111111;
    16'b0000100010000000: out_v[214] = 10'b1101000101;
    16'b0000100010001000: out_v[214] = 10'b1011011001;
    16'b0000101010001100: out_v[214] = 10'b1001001111;
    16'b0000111010011000: out_v[214] = 10'b0101111010;
    16'b0001101010001000: out_v[214] = 10'b0100110110;
    16'b0000100000001100: out_v[214] = 10'b1000100110;
    16'b0000000000001000: out_v[214] = 10'b1111000110;
    16'b0000111010011100: out_v[214] = 10'b0111011000;
    16'b0001111010001000: out_v[214] = 10'b1011101011;
    16'b0000001000001100: out_v[214] = 10'b0001001010;
    16'b0001111010011000: out_v[214] = 10'b1011101011;
    16'b0001111010011100: out_v[214] = 10'b1010011111;
    16'b0001111000000100: out_v[214] = 10'b1011110010;
    16'b0000011010011100: out_v[214] = 10'b1001111011;
    16'b0000111000001000: out_v[214] = 10'b0011100001;
    16'b0001001000001000: out_v[214] = 10'b1111111011;
    16'b0001101010011000: out_v[214] = 10'b0011011010;
    16'b0001101000011000: out_v[214] = 10'b0110101110;
    16'b0000101010010100: out_v[214] = 10'b0111000010;
    16'b0000100010010000: out_v[214] = 10'b1111100011;
    default: out_v[214] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000000001001: out_v[215] = 10'b0111000011;
    16'b0100001000001001: out_v[215] = 10'b1101010000;
    16'b0100011000011101: out_v[215] = 10'b0110101000;
    16'b0100010000001000: out_v[215] = 10'b0000010000;
    16'b0100001000011001: out_v[215] = 10'b0010011011;
    16'b0100001000011101: out_v[215] = 10'b1010011111;
    16'b0100000000011101: out_v[215] = 10'b0001000001;
    16'b0100010000000100: out_v[215] = 10'b1111110010;
    16'b0100000000001001: out_v[215] = 10'b1001000101;
    16'b0100000000011001: out_v[215] = 10'b0101110011;
    16'b0100010000001101: out_v[215] = 10'b0111001011;
    16'b0100000000001101: out_v[215] = 10'b0111011001;
    16'b0100010000001100: out_v[215] = 10'b1001100110;
    16'b0100010000011101: out_v[215] = 10'b0001000110;
    16'b0100011000011100: out_v[215] = 10'b1011100011;
    16'b0100001000000001: out_v[215] = 10'b1101000111;
    16'b0000001000000001: out_v[215] = 10'b1100011001;
    16'b0000001000001001: out_v[215] = 10'b0110100001;
    16'b0100000000001000: out_v[215] = 10'b0011010111;
    16'b0100001000010101: out_v[215] = 10'b0001110111;
    16'b0100011000001101: out_v[215] = 10'b0010011111;
    16'b0000010000011101: out_v[215] = 10'b1000101111;
    16'b0100010000011100: out_v[215] = 10'b1111101110;
    16'b0100001000010001: out_v[215] = 10'b1011110000;
    16'b0000011000011101: out_v[215] = 10'b1111010111;
    16'b0100000000001100: out_v[215] = 10'b1010010101;
    16'b0100001000001101: out_v[215] = 10'b1011001111;
    16'b0100010000001001: out_v[215] = 10'b0110000011;
    16'b0000000000011101: out_v[215] = 10'b1100011011;
    16'b0100011000001001: out_v[215] = 10'b0010001101;
    16'b0000010000010100: out_v[215] = 10'b1010111111;
    16'b0100011000001100: out_v[215] = 10'b0100011111;
    16'b0000000000001000: out_v[215] = 10'b1010100111;
    16'b0100010000000000: out_v[215] = 10'b1110010001;
    16'b0000010000011100: out_v[215] = 10'b0011110001;
    16'b0100011000001000: out_v[215] = 10'b0111111000;
    16'b0100001000011111: out_v[215] = 10'b0011001011;
    16'b0000001000000010: out_v[215] = 10'b0111000111;
    16'b0000001000000011: out_v[215] = 10'b0010010011;
    16'b0000001000001011: out_v[215] = 10'b1101010100;
    16'b0000000000000010: out_v[215] = 10'b1011001110;
    16'b0000000000000000: out_v[215] = 10'b0010011010;
    16'b0000000000000011: out_v[215] = 10'b1011011010;
    16'b0000000000001011: out_v[215] = 10'b0110111100;
    16'b0000011000001010: out_v[215] = 10'b1110100101;
    16'b0000011000000010: out_v[215] = 10'b0101100111;
    16'b0000011000001011: out_v[215] = 10'b0010000011;
    16'b0000001000000000: out_v[215] = 10'b0110001011;
    16'b0100001000000010: out_v[215] = 10'b0111100110;
    16'b0000001000010010: out_v[215] = 10'b0000100000;
    16'b0100001000011010: out_v[215] = 10'b0111100110;
    16'b0100001000010010: out_v[215] = 10'b1010100100;
    16'b0000001000001010: out_v[215] = 10'b1101000100;
    16'b0000010000001010: out_v[215] = 10'b1001001111;
    16'b0000011000011011: out_v[215] = 10'b0011001101;
    16'b0000001000011010: out_v[215] = 10'b0101000101;
    16'b0100001000001011: out_v[215] = 10'b0000110011;
    16'b0100000000010010: out_v[215] = 10'b1011100101;
    16'b0000011000001001: out_v[215] = 10'b1100011110;
    16'b0100011000000010: out_v[215] = 10'b1001010001;
    16'b0000011000001000: out_v[215] = 10'b1000000100;
    16'b0000011000011010: out_v[215] = 10'b0101010101;
    16'b0000001000011011: out_v[215] = 10'b1000101110;
    16'b0000000000010010: out_v[215] = 10'b0001101101;
    16'b0000000000011011: out_v[215] = 10'b1111101111;
    16'b0100001000001010: out_v[215] = 10'b0001011010;
    16'b0100001000011011: out_v[215] = 10'b1111110010;
    16'b0000010000001011: out_v[215] = 10'b0010001111;
    16'b0000001000001000: out_v[215] = 10'b1001011011;
    16'b0000010000000010: out_v[215] = 10'b0100110010;
    16'b0100000000000010: out_v[215] = 10'b1011101001;
    16'b0000000000001010: out_v[215] = 10'b1110010000;
    16'b0000011000000000: out_v[215] = 10'b1010100100;
    16'b0000010000001000: out_v[215] = 10'b1011011011;
    16'b0000000000000001: out_v[215] = 10'b0100001001;
    16'b0000001000010000: out_v[215] = 10'b0101011010;
    16'b0000010000001001: out_v[215] = 10'b0001110000;
    16'b0000010000000000: out_v[215] = 10'b1101110100;
    16'b0100000000000000: out_v[215] = 10'b0010011010;
    16'b0100000000000001: out_v[215] = 10'b1000100111;
    16'b0100010000001010: out_v[215] = 10'b1000101000;
    16'b0000001000011001: out_v[215] = 10'b0010110010;
    16'b0100010000001011: out_v[215] = 10'b1001101100;
    16'b0100001000000000: out_v[215] = 10'b0011100110;
    16'b0000001000010001: out_v[215] = 10'b0100101010;
    16'b0000001000011000: out_v[215] = 10'b1111000010;
    16'b0000000000010000: out_v[215] = 10'b1010101101;
    16'b0000010000000001: out_v[215] = 10'b1100001011;
    16'b0100010000000010: out_v[215] = 10'b0000111111;
    16'b0100010100000010: out_v[215] = 10'b1011001101;
    16'b0100011000001010: out_v[215] = 10'b0111011011;
    16'b0100000000001010: out_v[215] = 10'b1100011001;
    16'b0100011000000000: out_v[215] = 10'b1101011010;
    16'b0100000100000010: out_v[215] = 10'b0010110010;
    16'b0100011000001011: out_v[215] = 10'b0110000100;
    16'b0100001000000011: out_v[215] = 10'b0101010101;
    16'b0100000000001011: out_v[215] = 10'b1101010010;
    16'b0100001000001111: out_v[215] = 10'b0001011000;
    16'b0100001000001000: out_v[215] = 10'b0110010000;
    16'b0100000000000011: out_v[215] = 10'b1100110100;
    16'b0100011000000110: out_v[215] = 10'b0101000001;
    16'b0000000000011001: out_v[215] = 10'b1110111010;
    16'b0110001001001011: out_v[215] = 10'b1100001011;
    16'b0000001000010011: out_v[215] = 10'b1000111001;
    16'b0100001000001110: out_v[215] = 10'b1011000111;
    16'b0100011000001110: out_v[215] = 10'b0000011111;
    16'b0100011000000100: out_v[215] = 10'b0011111010;
    16'b0100011000001111: out_v[215] = 10'b1111000001;
    16'b0000011000001111: out_v[215] = 10'b0110001110;
    16'b0000010100001001: out_v[215] = 10'b0111100101;
    16'b0010001001001011: out_v[215] = 10'b0111010010;
    16'b0100010100001011: out_v[215] = 10'b1000100100;
    16'b0100010100001010: out_v[215] = 10'b1010101001;
    default: out_v[215] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100000000010100: out_v[216] = 10'b0000110110;
    16'b0000010101010100: out_v[216] = 10'b0110110111;
    16'b0101010101110100: out_v[216] = 10'b1001101111;
    16'b0101010101100100: out_v[216] = 10'b1101001000;
    16'b0100000100010100: out_v[216] = 10'b1000011011;
    16'b0000000101010100: out_v[216] = 10'b1000001011;
    16'b0101000101100100: out_v[216] = 10'b1111000101;
    16'b0001110101010100: out_v[216] = 10'b1110101101;
    16'b0101010101000100: out_v[216] = 10'b0101110001;
    16'b0100010100100100: out_v[216] = 10'b0001011011;
    16'b0100000101010100: out_v[216] = 10'b0110100110;
    16'b0001010101000100: out_v[216] = 10'b1100011011;
    16'b0100010101100100: out_v[216] = 10'b1000010011;
    16'b0100000100110100: out_v[216] = 10'b0011111101;
    16'b0101000100100100: out_v[216] = 10'b1001101110;
    16'b0001010101010100: out_v[216] = 10'b1011101110;
    16'b0000000100010100: out_v[216] = 10'b1011010011;
    16'b0101000101110100: out_v[216] = 10'b1000011111;
    16'b0000000101010000: out_v[216] = 10'b0000010000;
    16'b0101010001100100: out_v[216] = 10'b0111011011;
    16'b0100010100000100: out_v[216] = 10'b0110011011;
    16'b0000000101000100: out_v[216] = 10'b1111100010;
    16'b0100000100000100: out_v[216] = 10'b1111010001;
    16'b0000010101000100: out_v[216] = 10'b0011111011;
    16'b0000000100100100: out_v[216] = 10'b0001111011;
    16'b0100010101010100: out_v[216] = 10'b1100110110;
    16'b0100000101100100: out_v[216] = 10'b1110101011;
    16'b0001000101010100: out_v[216] = 10'b0011110111;
    16'b0000100101010100: out_v[216] = 10'b0100111100;
    16'b0100010101000100: out_v[216] = 10'b1010111111;
    16'b0101010000100100: out_v[216] = 10'b0100011011;
    16'b0101000101010100: out_v[216] = 10'b1011001110;
    16'b0100000100100100: out_v[216] = 10'b0100000001;
    16'b0101010101010100: out_v[216] = 10'b1000111111;
    16'b0101000101000100: out_v[216] = 10'b1110110101;
    16'b0000000001000100: out_v[216] = 10'b1101000101;
    16'b0101000000100100: out_v[216] = 10'b1000011001;
    16'b0100010101110100: out_v[216] = 10'b1110011001;
    16'b0100000101110100: out_v[216] = 10'b1010000001;
    16'b0000000001010100: out_v[216] = 10'b1000010010;
    16'b0101000001100100: out_v[216] = 10'b0110101001;
    16'b0001110100010100: out_v[216] = 10'b1111001011;
    16'b0101010100100100: out_v[216] = 10'b0011001110;
    16'b0100000101000100: out_v[216] = 10'b1110011111;
    16'b0000110101010100: out_v[216] = 10'b1000001110;
    16'b0000100000000100: out_v[216] = 10'b1010000101;
    16'b0000100001000000: out_v[216] = 10'b0110110111;
    16'b0000100000000000: out_v[216] = 10'b0100111001;
    16'b0000100001000100: out_v[216] = 10'b0100111000;
    16'b0000000000000100: out_v[216] = 10'b1100011011;
    16'b0100100001000000: out_v[216] = 10'b1000100011;
    16'b0000000000000000: out_v[216] = 10'b1011000010;
    16'b0100100001000100: out_v[216] = 10'b1011010101;
    16'b0100100000000000: out_v[216] = 10'b1001010111;
    16'b0100100000000100: out_v[216] = 10'b1100111010;
    16'b0100100000100100: out_v[216] = 10'b0010111000;
    16'b0000100001010100: out_v[216] = 10'b1011000010;
    16'b0100100001100000: out_v[216] = 10'b1100000101;
    16'b0100100001100100: out_v[216] = 10'b0010010110;
    16'b0100100100000100: out_v[216] = 10'b0010111111;
    16'b0000100100000100: out_v[216] = 10'b1001001001;
    16'b0000100000010100: out_v[216] = 10'b0011001100;
    16'b0100000001000100: out_v[216] = 10'b0010001100;
    16'b0101110100010100: out_v[216] = 10'b1011100100;
    16'b0101100101000100: out_v[216] = 10'b0111011100;
    16'b0101100101010100: out_v[216] = 10'b1000010010;
    16'b0101100100000100: out_v[216] = 10'b0101110111;
    16'b0000100100010100: out_v[216] = 10'b0001110011;
    16'b0000100000100100: out_v[216] = 10'b0001110111;
    16'b0100100101000100: out_v[216] = 10'b1000011110;
    16'b0001100100000100: out_v[216] = 10'b1101010111;
    16'b0100100001110100: out_v[216] = 10'b1100110111;
    16'b0000100001110100: out_v[216] = 10'b0111001010;
    16'b0100100001010100: out_v[216] = 10'b0000101110;
    16'b0100000001100100: out_v[216] = 10'b1011110010;
    16'b0001100100010100: out_v[216] = 10'b0111110111;
    16'b0100000001000000: out_v[216] = 10'b0000111100;
    16'b0100100100010100: out_v[216] = 10'b1100010000;
    16'b0100100100000000: out_v[216] = 10'b0101011010;
    16'b0000100000100000: out_v[216] = 10'b1001000101;
    16'b0100000000000100: out_v[216] = 10'b0111000111;
    16'b0000100101000100: out_v[216] = 10'b1110010110;
    16'b0000100100010000: out_v[216] = 10'b1101000111;
    16'b0000100100000000: out_v[216] = 10'b0011010100;
    16'b0000100000010000: out_v[216] = 10'b0011000101;
    16'b0100100101010100: out_v[216] = 10'b0011001111;
    16'b0000100001100100: out_v[216] = 10'b0111101001;
    16'b0000100000110100: out_v[216] = 10'b0111100101;
    16'b0100100101100100: out_v[216] = 10'b0111100100;
    16'b0100000000110100: out_v[216] = 10'b1001011011;
    16'b0100000001010100: out_v[216] = 10'b0111000100;
    16'b0000000001000000: out_v[216] = 10'b1001011001;
    16'b0100000000100100: out_v[216] = 10'b0111100000;
    16'b0000000001010000: out_v[216] = 10'b0111011000;
    16'b0100000000010000: out_v[216] = 10'b1001100101;
    16'b0100000000000000: out_v[216] = 10'b0111011010;
    16'b0100000001010000: out_v[216] = 10'b1001110000;
    16'b0100000001110100: out_v[216] = 10'b1101011010;
    16'b0100000100010000: out_v[216] = 10'b0011011111;
    16'b0000000001110100: out_v[216] = 10'b0111011110;
    16'b0000000000010100: out_v[216] = 10'b0001111001;
    16'b0100000000110000: out_v[216] = 10'b1010100111;
    16'b0000100100110100: out_v[216] = 10'b0110111001;
    16'b0000100100100100: out_v[216] = 10'b1100000101;
    16'b0000100101000000: out_v[216] = 10'b0110111110;
    16'b0000110101010000: out_v[216] = 10'b0001010001;
    16'b0101100100110100: out_v[216] = 10'b1001001111;
    16'b0000100100110000: out_v[216] = 10'b1011001110;
    16'b0000100101100000: out_v[216] = 10'b1010101101;
    16'b0000100101010000: out_v[216] = 10'b0001110000;
    16'b0100100100110000: out_v[216] = 10'b1000011011;
    16'b0001100101000000: out_v[216] = 10'b1111001010;
    16'b0001100100010000: out_v[216] = 10'b0100001111;
    16'b0000100101100100: out_v[216] = 10'b0000011011;
    16'b0100000100110000: out_v[216] = 10'b1000110111;
    16'b0000110100000000: out_v[216] = 10'b0010111011;
    16'b0000000101100000: out_v[216] = 10'b0001110011;
    16'b0000100101110000: out_v[216] = 10'b0111101100;
    16'b0101100100110000: out_v[216] = 10'b0110111111;
    16'b0100100100110100: out_v[216] = 10'b1000111111;
    16'b0000100101110100: out_v[216] = 10'b1001010010;
    16'b0001110101010000: out_v[216] = 10'b1111101110;
    16'b0001110100010000: out_v[216] = 10'b1000111011;
    16'b0101000100110100: out_v[216] = 10'b0001110111;
    16'b0000110100010000: out_v[216] = 10'b1010010100;
    16'b0001100101110000: out_v[216] = 10'b0110101111;
    16'b0000000101000000: out_v[216] = 10'b0111110000;
    16'b0001100101010100: out_v[216] = 10'b0101010110;
    16'b0000000101100100: out_v[216] = 10'b0000111011;
    16'b0001100101010000: out_v[216] = 10'b0110101100;
    16'b0000000100000100: out_v[216] = 10'b0001111011;
    16'b0001110101110000: out_v[216] = 10'b1010111001;
    16'b0000110101110000: out_v[216] = 10'b0010111101;
    16'b0100100100010000: out_v[216] = 10'b0110011001;
    16'b0001100100000000: out_v[216] = 10'b0111100110;
    16'b0000110001000100: out_v[216] = 10'b0111111100;
    16'b0000110101000100: out_v[216] = 10'b1011100010;
    16'b0100000001110000: out_v[216] = 10'b1010101001;
    16'b0100000000100000: out_v[216] = 10'b0001110001;
    16'b0000110001000000: out_v[216] = 10'b0010001111;
    16'b0000110000000000: out_v[216] = 10'b0011001101;
    16'b0000000001100100: out_v[216] = 10'b0101110110;
    16'b0000110101000000: out_v[216] = 10'b0100001011;
    16'b0100100100100100: out_v[216] = 10'b1100101011;
    16'b0000010001000100: out_v[216] = 10'b1011010011;
    16'b0100100101010000: out_v[216] = 10'b0101001001;
    16'b0100100101000000: out_v[216] = 10'b0011010111;
    16'b0100100101110000: out_v[216] = 10'b1001001000;
    16'b0100100001010000: out_v[216] = 10'b0111101101;
    16'b0100100101100000: out_v[216] = 10'b0111011000;
    16'b0100000101100000: out_v[216] = 10'b0001100000;
    16'b0000100001010000: out_v[216] = 10'b1001001011;
    16'b0100000101010000: out_v[216] = 10'b1101110110;
    16'b0100000101000000: out_v[216] = 10'b0001010101;
    16'b0100000101110000: out_v[216] = 10'b1001001011;
    16'b0000110001110100: out_v[216] = 10'b0111001001;
    16'b0000100001110000: out_v[216] = 10'b1000000111;
    16'b0000000001110000: out_v[216] = 10'b0110001100;
    16'b0000100001100000: out_v[216] = 10'b1110100000;
    16'b0000000001100000: out_v[216] = 10'b1000010111;
    16'b0000110000100100: out_v[216] = 10'b1001100110;
    16'b0000000000110000: out_v[216] = 10'b1100100111;
    16'b0000110000000100: out_v[216] = 10'b1101000100;
    16'b0000110000100000: out_v[216] = 10'b0011010110;
    16'b0000110001110000: out_v[216] = 10'b1011011100;
    16'b0000110000110100: out_v[216] = 10'b0100011110;
    16'b0000110100000100: out_v[216] = 10'b1111100000;
    16'b0000110001100100: out_v[216] = 10'b0110100011;
    16'b0100110000100100: out_v[216] = 10'b1101011111;
    16'b0100100000100000: out_v[216] = 10'b0100001010;
    16'b0000110101100100: out_v[216] = 10'b0111100011;
    16'b0100100000110100: out_v[216] = 10'b0101001010;
    16'b0000000000100100: out_v[216] = 10'b0101011000;
    16'b0000000101110100: out_v[216] = 10'b1100100010;
    16'b0100100100110110: out_v[216] = 10'b1001101101;
    16'b0100100100110010: out_v[216] = 10'b1011101111;
    default: out_v[216] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010000000001000: out_v[217] = 10'b0111010101;
    16'b0001100000000100: out_v[217] = 10'b1000010011;
    16'b0001100001001100: out_v[217] = 10'b1111011110;
    16'b0011100000001100: out_v[217] = 10'b1000001100;
    16'b0010000000001100: out_v[217] = 10'b0100111010;
    16'b0001000000000000: out_v[217] = 10'b0111010011;
    16'b0001100000001000: out_v[217] = 10'b0100111011;
    16'b0001000000000100: out_v[217] = 10'b1111111010;
    16'b0001100000000000: out_v[217] = 10'b1100010111;
    16'b0011100001001000: out_v[217] = 10'b0010111111;
    16'b0000100000000100: out_v[217] = 10'b1010011011;
    16'b0011100000000100: out_v[217] = 10'b0100101101;
    16'b0001100001000100: out_v[217] = 10'b1000000011;
    16'b0001100000001100: out_v[217] = 10'b1000001111;
    16'b0011000000001100: out_v[217] = 10'b0110101010;
    16'b0011100001000100: out_v[217] = 10'b1100010110;
    16'b0001000000001000: out_v[217] = 10'b0011000100;
    16'b0011100001001100: out_v[217] = 10'b1000000001;
    16'b0011000000000100: out_v[217] = 10'b0111001011;
    16'b1001000000000000: out_v[217] = 10'b1011100111;
    16'b0011000000000000: out_v[217] = 10'b1100100111;
    16'b0000000000000000: out_v[217] = 10'b1110110110;
    16'b0001100001000000: out_v[217] = 10'b0001111111;
    16'b0011100000001000: out_v[217] = 10'b1111101010;
    16'b0011000000001000: out_v[217] = 10'b1011011100;
    16'b0000100001001100: out_v[217] = 10'b1110001010;
    16'b0000100001000100: out_v[217] = 10'b1010011111;
    16'b0011000001001000: out_v[217] = 10'b1100011011;
    16'b0010100000001100: out_v[217] = 10'b1000000111;
    16'b0001100001001000: out_v[217] = 10'b0010101101;
    16'b0010000000000000: out_v[217] = 10'b1110110000;
    16'b0000100000001100: out_v[217] = 10'b0010100110;
    16'b1011000000000000: out_v[217] = 10'b1110001100;
    16'b0001000000001100: out_v[217] = 10'b0011110001;
    16'b0001000001001000: out_v[217] = 10'b1001010011;
    16'b1001100001000100: out_v[217] = 10'b0101101101;
    16'b1000000000000000: out_v[217] = 10'b1010110011;
    16'b0000000000001000: out_v[217] = 10'b0100111100;
    16'b1010000000000000: out_v[217] = 10'b1110001101;
    16'b1010000000001000: out_v[217] = 10'b1100000110;
    16'b1000000000001000: out_v[217] = 10'b0000011111;
    16'b1111000000001000: out_v[217] = 10'b1111110100;
    16'b1011000000010000: out_v[217] = 10'b1110100011;
    16'b0111000000000000: out_v[217] = 10'b1010111110;
    16'b1111000000010000: out_v[217] = 10'b1111110010;
    16'b1101000000010000: out_v[217] = 10'b0110100101;
    16'b1011000000011000: out_v[217] = 10'b0111110011;
    16'b1011000000001000: out_v[217] = 10'b1100010000;
    16'b1111000000000000: out_v[217] = 10'b1010001110;
    16'b1001000000000100: out_v[217] = 10'b0111110100;
    16'b0011000000011000: out_v[217] = 10'b1010000111;
    16'b0111000000010000: out_v[217] = 10'b0100111011;
    16'b1010000000010000: out_v[217] = 10'b1110100000;
    16'b1001000000010000: out_v[217] = 10'b0011001011;
    16'b1001000000001000: out_v[217] = 10'b1011001110;
    16'b0111000000001000: out_v[217] = 10'b0000011111;
    16'b1111000000000100: out_v[217] = 10'b0111101010;
    16'b0111000000011000: out_v[217] = 10'b0010011010;
    16'b1011100000000100: out_v[217] = 10'b1001000110;
    16'b0011000000010000: out_v[217] = 10'b1010110011;
    16'b1000000000000100: out_v[217] = 10'b0110010100;
    16'b1011000000000100: out_v[217] = 10'b1100011110;
    16'b1111000000011000: out_v[217] = 10'b1110000111;
    16'b1010000000001100: out_v[217] = 10'b1000111000;
    16'b1000000000001100: out_v[217] = 10'b1010101010;
    16'b1011000000001100: out_v[217] = 10'b0111001011;
    16'b0000000000001100: out_v[217] = 10'b0001101001;
    16'b0010000000000100: out_v[217] = 10'b1101001001;
    16'b1010000000000100: out_v[217] = 10'b0011111000;
    16'b1000100000000100: out_v[217] = 10'b0010010010;
    16'b1001000000001100: out_v[217] = 10'b0011110010;
    16'b1000100000001100: out_v[217] = 10'b1001000110;
    16'b1000100000001000: out_v[217] = 10'b0000110111;
    16'b1000100000000000: out_v[217] = 10'b0010010010;
    16'b0001000001000000: out_v[217] = 10'b1000111011;
    16'b0010000000011000: out_v[217] = 10'b0001000010;
    16'b1001000000010100: out_v[217] = 10'b1011101111;
    16'b1100100000000100: out_v[217] = 10'b1101101111;
    16'b1011100000010100: out_v[217] = 10'b1011010100;
    16'b1010000000011000: out_v[217] = 10'b1100100010;
    16'b1011000000010100: out_v[217] = 10'b1011100101;
    16'b1010000000010100: out_v[217] = 10'b1000111001;
    16'b0010000000010000: out_v[217] = 10'b1001000110;
    16'b0010000000010100: out_v[217] = 10'b1100111010;
    16'b0011100000010100: out_v[217] = 10'b0111110110;
    16'b1011000000011100: out_v[217] = 10'b1011011010;
    16'b1000000000010000: out_v[217] = 10'b0111101100;
    16'b0010000000011100: out_v[217] = 10'b1111011011;
    16'b1010000000011100: out_v[217] = 10'b1011111100;
    16'b0100000000000100: out_v[217] = 10'b0111110001;
    16'b0011000000010100: out_v[217] = 10'b1011111011;
    16'b1001100000000100: out_v[217] = 10'b1111000110;
    16'b1111100000000100: out_v[217] = 10'b1101111011;
    16'b1101100000000100: out_v[217] = 10'b1011100001;
    16'b0000000000010000: out_v[217] = 10'b1011011011;
    16'b1110000000000100: out_v[217] = 10'b0111101111;
    16'b1100000000000100: out_v[217] = 10'b1101101010;
    16'b1000000100001001: out_v[217] = 10'b0010011111;
    16'b0000000100001001: out_v[217] = 10'b1111011011;
    16'b1000000000000001: out_v[217] = 10'b1101000100;
    16'b1000000100000001: out_v[217] = 10'b1001101100;
    16'b1001000001000000: out_v[217] = 10'b0001110110;
    16'b1001100001000000: out_v[217] = 10'b0110000111;
    default: out_v[217] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100111000000000: out_v[218] = 10'b0000011101;
    16'b0000001000001000: out_v[218] = 10'b0110100011;
    16'b0100001000001000: out_v[218] = 10'b1010000001;
    16'b0110010000001000: out_v[218] = 10'b0011001011;
    16'b0110111000000000: out_v[218] = 10'b0111000101;
    16'b0000001000000000: out_v[218] = 10'b1111100001;
    16'b0100011001000000: out_v[218] = 10'b0010111101;
    16'b0100001001000000: out_v[218] = 10'b0000000101;
    16'b0110010001001000: out_v[218] = 10'b1011001001;
    16'b0010111000000000: out_v[218] = 10'b0011110011;
    16'b0100101000001000: out_v[218] = 10'b1000111011;
    16'b0100001000000000: out_v[218] = 10'b1010000010;
    16'b0100011000001000: out_v[218] = 10'b0100110100;
    16'b0100101000000000: out_v[218] = 10'b1001000011;
    16'b0000011000000000: out_v[218] = 10'b1100111000;
    16'b0100010000000000: out_v[218] = 10'b1110001100;
    16'b0110010000000000: out_v[218] = 10'b0001011010;
    16'b0100010000001000: out_v[218] = 10'b1100111011;
    16'b0010011000001000: out_v[218] = 10'b1111111010;
    16'b0100011000000000: out_v[218] = 10'b0100010100;
    16'b0000011000001000: out_v[218] = 10'b1000111101;
    16'b0100011001001000: out_v[218] = 10'b0100101011;
    16'b0000111000000000: out_v[218] = 10'b0100011110;
    16'b0110011001000000: out_v[218] = 10'b1001110110;
    16'b0100010001000000: out_v[218] = 10'b0010100101;
    16'b0100010001001000: out_v[218] = 10'b1000011101;
    16'b0000010001000000: out_v[218] = 10'b0000000111;
    16'b0000010001001000: out_v[218] = 10'b1111011001;
    16'b0000101000000000: out_v[218] = 10'b1001000001;
    16'b0110011000001000: out_v[218] = 10'b0101110110;
    16'b0010010001000000: out_v[218] = 10'b1011111000;
    16'b0110010001000000: out_v[218] = 10'b0111000010;
    16'b0000010000000000: out_v[218] = 10'b1010001101;
    16'b0100111001001000: out_v[218] = 10'b0101011011;
    16'b0000010000001000: out_v[218] = 10'b0010000110;
    16'b0000111000001000: out_v[218] = 10'b0100010110;
    16'b0110011001001000: out_v[218] = 10'b1011100011;
    16'b0010010000000000: out_v[218] = 10'b0101110101;
    16'b0010011000000000: out_v[218] = 10'b0111111000;
    16'b0000101000001000: out_v[218] = 10'b1111101001;
    16'b0110011000000000: out_v[218] = 10'b1010111010;
    16'b0100001001001000: out_v[218] = 10'b1011100111;
    16'b0100111000001000: out_v[218] = 10'b1001100010;
    16'b0110111000001000: out_v[218] = 10'b1111010001;
    16'b0000100000000000: out_v[218] = 10'b0110110010;
    16'b0000000000000000: out_v[218] = 10'b0111111011;
    16'b0010000000000000: out_v[218] = 10'b1001100100;
    16'b0000100000001000: out_v[218] = 10'b1000000100;
    16'b0110110000000000: out_v[218] = 10'b0111000110;
    16'b0010110000000000: out_v[218] = 10'b0111000100;
    16'b0110110001000000: out_v[218] = 10'b1011110001;
    16'b0000110000000000: out_v[218] = 10'b1011001100;
    16'b0100110001000000: out_v[218] = 10'b0001110111;
    16'b0110000000000000: out_v[218] = 10'b1111011011;
    16'b0000100001000000: out_v[218] = 10'b0000111010;
    16'b0010100000000000: out_v[218] = 10'b0010110110;
    16'b0010010000001000: out_v[218] = 10'b0001100001;
    16'b0110100000000000: out_v[218] = 10'b1010100101;
    16'b0110110000001000: out_v[218] = 10'b1000011111;
    16'b0100110000000000: out_v[218] = 10'b0100101100;
    16'b0010110001000000: out_v[218] = 10'b0111101000;
    16'b0000110001000000: out_v[218] = 10'b0110110010;
    16'b0010110000001000: out_v[218] = 10'b1011110110;
    16'b0100110000001000: out_v[218] = 10'b1101101100;
    16'b0000110000001000: out_v[218] = 10'b0100111100;
    16'b0000101001000000: out_v[218] = 10'b0000011110;
    16'b0110100000001000: out_v[218] = 10'b1011011110;
    16'b0110111001000000: out_v[218] = 10'b1101110000;
    16'b0100111001000000: out_v[218] = 10'b0010001111;
    16'b0000111001000000: out_v[218] = 10'b0111001110;
    16'b0000011001000000: out_v[218] = 10'b1110111000;
    16'b0110001000000000: out_v[218] = 10'b0100001100;
    16'b0010001000000000: out_v[218] = 10'b1010011000;
    16'b0100100000000000: out_v[218] = 10'b0000111001;
    16'b0100100000001000: out_v[218] = 10'b0001011100;
    16'b0100000000001000: out_v[218] = 10'b0011111110;
    16'b0000000000001000: out_v[218] = 10'b0110110000;
    16'b0100000000000000: out_v[218] = 10'b0111110010;
    16'b0100100001000000: out_v[218] = 10'b0011111010;
    16'b0100000001000000: out_v[218] = 10'b1001000011;
    16'b0000000000001001: out_v[218] = 10'b0111011011;
    16'b0000001000001001: out_v[218] = 10'b0011001010;
    16'b0000000000000001: out_v[218] = 10'b0111011101;
    16'b0000010000000001: out_v[218] = 10'b0111110000;
    16'b0010111000001000: out_v[218] = 10'b1111000011;
    16'b0100110010000000: out_v[218] = 10'b1011000111;
    default: out_v[218] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000100010000000: out_v[219] = 10'b0000101101;
    16'b0000100011010000: out_v[219] = 10'b0011001110;
    16'b1000100111010000: out_v[219] = 10'b0000010001;
    16'b1000100111000000: out_v[219] = 10'b0110011000;
    16'b0000100111010000: out_v[219] = 10'b1101001001;
    16'b0000100111000000: out_v[219] = 10'b0000000011;
    16'b0000000010010000: out_v[219] = 10'b1010010111;
    16'b0000000011000000: out_v[219] = 10'b1011100100;
    16'b0000100101000000: out_v[219] = 10'b1001000011;
    16'b0000100111110000: out_v[219] = 10'b1111100101;
    16'b0000100010010000: out_v[219] = 10'b0111001001;
    16'b1000000101000000: out_v[219] = 10'b0011010011;
    16'b1000100101000000: out_v[219] = 10'b0010101000;
    16'b0000100011000000: out_v[219] = 10'b0010010101;
    16'b0000000011010000: out_v[219] = 10'b0010110110;
    16'b0000100100000000: out_v[219] = 10'b1011011011;
    16'b0000100110000000: out_v[219] = 10'b1101110100;
    16'b1000100100000000: out_v[219] = 10'b1010000110;
    16'b0000000011110000: out_v[219] = 10'b0011101010;
    16'b1000000111000000: out_v[219] = 10'b0110100101;
    16'b1000100110000000: out_v[219] = 10'b0010001011;
    16'b0000100101010000: out_v[219] = 10'b1011011011;
    16'b0000100110010000: out_v[219] = 10'b0010011100;
    16'b0000100000000000: out_v[219] = 10'b0011110001;
    16'b0000000001010000: out_v[219] = 10'b1000011101;
    16'b0000000010000000: out_v[219] = 10'b0001011001;
    16'b1000100110010000: out_v[219] = 10'b0010011100;
    16'b0000100001000000: out_v[219] = 10'b0111100000;
    16'b0100000000100000: out_v[219] = 10'b1000010011;
    16'b0100000010100000: out_v[219] = 10'b1100011011;
    16'b0100000010110000: out_v[219] = 10'b0101011010;
    16'b0100000001100000: out_v[219] = 10'b1100011000;
    16'b0100000000110000: out_v[219] = 10'b1101100110;
    16'b0100000001000000: out_v[219] = 10'b0100010100;
    16'b0100000000000000: out_v[219] = 10'b1110011101;
    16'b0100100010110000: out_v[219] = 10'b0001000010;
    16'b0100000011010000: out_v[219] = 10'b1011011010;
    16'b0100000010010000: out_v[219] = 10'b1110111000;
    16'b0100000010000000: out_v[219] = 10'b1001000100;
    16'b0100000011100000: out_v[219] = 10'b1011101001;
    16'b0100000001010000: out_v[219] = 10'b0001110100;
    16'b0100000011110000: out_v[219] = 10'b1111011000;
    16'b0000000000010000: out_v[219] = 10'b0010001100;
    16'b0100000001110000: out_v[219] = 10'b0111001001;
    16'b0100000000010000: out_v[219] = 10'b1011001001;
    16'b0100000011000000: out_v[219] = 10'b0001000100;
    16'b0100100001010000: out_v[219] = 10'b0011101111;
    16'b0000000001000000: out_v[219] = 10'b1101001100;
    16'b0000100001010000: out_v[219] = 10'b1101101110;
    16'b0100100011010000: out_v[219] = 10'b1000111111;
    16'b0000000000000000: out_v[219] = 10'b0010111100;
    16'b0000100011110000: out_v[219] = 10'b0000101110;
    16'b0000000010100000: out_v[219] = 10'b1101111100;
    16'b0101000010110000: out_v[219] = 10'b0101011111;
    16'b0100100010100000: out_v[219] = 10'b1100000000;
    16'b0100100011110000: out_v[219] = 10'b1100101111;
    16'b0000100011100000: out_v[219] = 10'b0011111001;
    16'b0100100011100000: out_v[219] = 10'b0100011010;
    16'b0000000010110000: out_v[219] = 10'b1001101100;
    16'b0000000001100000: out_v[219] = 10'b1010111000;
    16'b0000000011100000: out_v[219] = 10'b0110100010;
    16'b0000000000100000: out_v[219] = 10'b1101110001;
    16'b0100100000100000: out_v[219] = 10'b1001011001;
    16'b0101000010100000: out_v[219] = 10'b0101110010;
    16'b0101000010010000: out_v[219] = 10'b0001011100;
    16'b0100100110010000: out_v[219] = 10'b1100001001;
    16'b0100100100010000: out_v[219] = 10'b1001001011;
    16'b0100100100000000: out_v[219] = 10'b0000111110;
    16'b1000100100010000: out_v[219] = 10'b1101111010;
    16'b0100100000010000: out_v[219] = 10'b1111011101;
    16'b0100100000000000: out_v[219] = 10'b1011110000;
    16'b1100100110010000: out_v[219] = 10'b0100001110;
    16'b1100100100010000: out_v[219] = 10'b1001110110;
    16'b0100100010010000: out_v[219] = 10'b1101000100;
    16'b1100100100000000: out_v[219] = 10'b0110111110;
    16'b0000100000010000: out_v[219] = 10'b0110111010;
    16'b1000000100000000: out_v[219] = 10'b0011011011;
    16'b1000000110010000: out_v[219] = 10'b1101001011;
    16'b1100100110110000: out_v[219] = 10'b0101010111;
    16'b1100000100000000: out_v[219] = 10'b1100110001;
    16'b0100100110110000: out_v[219] = 10'b1100000111;
    16'b1100000110010000: out_v[219] = 10'b1101100010;
    16'b1000000100010000: out_v[219] = 10'b1000010010;
    16'b0000100100010000: out_v[219] = 10'b0110111011;
    16'b0100100010000000: out_v[219] = 10'b0011001011;
    16'b0100100110000000: out_v[219] = 10'b1100111101;
    16'b0100100111010000: out_v[219] = 10'b1101000100;
    16'b0100100011000000: out_v[219] = 10'b0010011001;
    16'b0000100100100000: out_v[219] = 10'b1001001000;
    16'b0100100001100000: out_v[219] = 10'b1101000011;
    16'b0100100001000000: out_v[219] = 10'b0101111010;
    16'b0100100111110000: out_v[219] = 10'b0011111110;
    16'b0000100010100000: out_v[219] = 10'b0011110110;
    16'b0000100000100000: out_v[219] = 10'b0011100110;
    16'b0000100001100000: out_v[219] = 10'b1111100110;
    16'b0000100010110000: out_v[219] = 10'b1000100000;
    16'b0100101010000000: out_v[219] = 10'b1111111010;
    16'b0100001010010000: out_v[219] = 10'b1101000100;
    16'b0000101010010000: out_v[219] = 10'b1111100111;
    16'b0100101010010000: out_v[219] = 10'b1000011111;
    16'b0000001010010000: out_v[219] = 10'b0111101101;
    16'b0100101110010000: out_v[219] = 10'b1110100111;
    16'b0100101111010000: out_v[219] = 10'b1101101001;
    16'b0100100111000000: out_v[219] = 10'b1011010111;
    16'b0000101110010000: out_v[219] = 10'b1111100110;
    16'b1100100111010000: out_v[219] = 10'b0111110101;
    16'b0100001010000000: out_v[219] = 10'b0101111110;
    16'b0100101010110000: out_v[219] = 10'b1001011100;
    16'b1000100000010000: out_v[219] = 10'b0111000111;
    16'b1000100110110000: out_v[219] = 10'b1110100011;
    16'b1000100010010000: out_v[219] = 10'b0100110010;
    16'b1000000010010000: out_v[219] = 10'b0011110010;
    16'b1100100010010000: out_v[219] = 10'b1101010100;
    16'b1000000000010000: out_v[219] = 10'b1001001010;
    16'b1000100000000000: out_v[219] = 10'b1100100010;
    16'b1000100010110000: out_v[219] = 10'b1111000100;
    16'b1100100000010000: out_v[219] = 10'b0111001111;
    16'b0100100000110000: out_v[219] = 10'b1100010001;
    16'b1100100000100000: out_v[219] = 10'b0111000010;
    default: out_v[219] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1000100000100010: out_v[220] = 10'b0010110111;
    16'b1100100000100000: out_v[220] = 10'b1110011111;
    16'b1000100000100000: out_v[220] = 10'b0100010011;
    16'b0000100000100010: out_v[220] = 10'b0010100111;
    16'b1100100000000010: out_v[220] = 10'b1110000001;
    16'b1100000000000000: out_v[220] = 10'b1101110000;
    16'b0000100000000010: out_v[220] = 10'b1110110000;
    16'b1000000100100000: out_v[220] = 10'b0110111011;
    16'b1100000000100010: out_v[220] = 10'b1100001011;
    16'b0000000000100010: out_v[220] = 10'b1100000101;
    16'b1100000000000010: out_v[220] = 10'b1011110010;
    16'b1010100000100010: out_v[220] = 10'b0101011001;
    16'b1100100000100010: out_v[220] = 10'b0110010011;
    16'b1000100100100000: out_v[220] = 10'b0010111011;
    16'b1000000000100010: out_v[220] = 10'b0011100011;
    16'b0000100100100010: out_v[220] = 10'b0101110110;
    16'b1000100100100010: out_v[220] = 10'b0101011101;
    16'b1000000000100000: out_v[220] = 10'b1011010111;
    16'b0100100000000010: out_v[220] = 10'b1001111011;
    16'b1100000000100000: out_v[220] = 10'b1010111000;
    16'b0000100000000000: out_v[220] = 10'b1010100011;
    16'b0000100110100000: out_v[220] = 10'b1010011011;
    16'b0000100100100000: out_v[220] = 10'b0110110011;
    16'b1000100010100010: out_v[220] = 10'b1111000101;
    16'b1000100110100000: out_v[220] = 10'b1011011001;
    16'b0100100000100010: out_v[220] = 10'b1001001001;
    16'b1100100000000000: out_v[220] = 10'b0111001111;
    16'b1000100010100000: out_v[220] = 10'b1111000111;
    16'b0000100000100000: out_v[220] = 10'b1110011001;
    16'b1100100100100010: out_v[220] = 10'b1011011011;
    16'b1000100000000000: out_v[220] = 10'b1110010011;
    16'b1100100100100000: out_v[220] = 10'b0101110110;
    16'b1000100110100010: out_v[220] = 10'b0010011101;
    16'b0000100110100010: out_v[220] = 10'b0101110011;
    16'b1110100000100010: out_v[220] = 10'b0000010001;
    16'b1010101000000010: out_v[220] = 10'b0101010110;
    16'b0010001000000010: out_v[220] = 10'b0100010100;
    16'b0000001000000010: out_v[220] = 10'b0000110010;
    16'b1000101000000010: out_v[220] = 10'b0001000100;
    16'b0010000000000010: out_v[220] = 10'b1110001001;
    16'b1010101000000000: out_v[220] = 10'b1100011101;
    16'b0000001000000000: out_v[220] = 10'b0001000010;
    16'b1000101000000000: out_v[220] = 10'b1110101101;
    16'b0010101000000010: out_v[220] = 10'b1110110001;
    16'b1000001000000010: out_v[220] = 10'b0111000011;
    16'b0010101000000000: out_v[220] = 10'b0100011010;
    16'b0000000000000010: out_v[220] = 10'b0010001010;
    16'b1010101000100010: out_v[220] = 10'b1001101110;
    16'b1010001000000010: out_v[220] = 10'b1101000001;
    16'b0010001000000000: out_v[220] = 10'b0111010001;
    16'b1010100000100000: out_v[220] = 10'b1101011110;
    16'b0010101100000000: out_v[220] = 10'b1000001101;
    16'b1010101100000010: out_v[220] = 10'b1001100001;
    16'b1010101000100000: out_v[220] = 10'b1010101111;
    16'b0010001110000010: out_v[220] = 10'b1110100101;
    16'b1110101000000000: out_v[220] = 10'b0111110001;
    16'b0000001100000010: out_v[220] = 10'b1110011001;
    16'b1110101000100010: out_v[220] = 10'b1101001100;
    16'b0010101100100000: out_v[220] = 10'b0000011111;
    16'b1010101110100000: out_v[220] = 10'b1110100010;
    16'b1100101000100000: out_v[220] = 10'b0000101110;
    16'b0010101000100010: out_v[220] = 10'b1001001010;
    16'b1110101000100000: out_v[220] = 10'b1100100111;
    16'b1110101100100000: out_v[220] = 10'b1011110101;
    16'b1000101100100000: out_v[220] = 10'b1100011110;
    16'b0010001000100010: out_v[220] = 10'b0001011100;
    16'b1010101100100000: out_v[220] = 10'b0010100011;
    16'b1110101010100000: out_v[220] = 10'b0111111011;
    16'b0000001000100010: out_v[220] = 10'b0101010101;
    16'b0010101000100000: out_v[220] = 10'b0001101010;
    16'b1010101100000000: out_v[220] = 10'b0101011001;
    16'b1010101110000000: out_v[220] = 10'b0101000011;
    16'b1010101010000000: out_v[220] = 10'b0011111101;
    16'b0010101100100010: out_v[220] = 10'b0111101010;
    16'b1110001000100000: out_v[220] = 10'b0101000101;
    16'b0110001000100000: out_v[220] = 10'b1110110011;
    16'b0010001100000010: out_v[220] = 10'b0100111111;
    16'b1110101110100000: out_v[220] = 10'b1101010011;
    16'b1110101010100010: out_v[220] = 10'b0010011100;
    16'b1100101100100000: out_v[220] = 10'b1001101111;
    16'b1110101100100010: out_v[220] = 10'b0111011111;
    16'b0010001100100010: out_v[220] = 10'b1011000010;
    16'b1010101110000010: out_v[220] = 10'b0001011111;
    16'b0010101100000010: out_v[220] = 10'b0010100100;
    16'b1000101000100000: out_v[220] = 10'b0001110010;
    16'b1010101010100000: out_v[220] = 10'b0011001101;
    16'b0000001100100010: out_v[220] = 10'b1001000110;
    16'b1100001000100000: out_v[220] = 10'b0001010110;
    16'b1010101100100010: out_v[220] = 10'b0110111010;
    16'b0010101110000010: out_v[220] = 10'b0101100000;
    16'b1010100100000010: out_v[220] = 10'b0000011011;
    16'b1110100000000010: out_v[220] = 10'b0000010001;
    16'b0010000010000010: out_v[220] = 10'b0010010111;
    16'b1110100100000000: out_v[220] = 10'b1110110011;
    16'b1110000000000000: out_v[220] = 10'b1010011100;
    16'b1010100110000000: out_v[220] = 10'b0011111011;
    16'b1010100100000000: out_v[220] = 10'b0010110110;
    16'b0010000100000010: out_v[220] = 10'b0110011101;
    16'b1010100000000000: out_v[220] = 10'b1000011110;
    16'b1110100000000000: out_v[220] = 10'b0011001011;
    16'b0010000110000010: out_v[220] = 10'b0011011111;
    16'b0010100100000010: out_v[220] = 10'b1100110111;
    16'b1110101000000010: out_v[220] = 10'b1010001110;
    16'b1010100000000010: out_v[220] = 10'b1001011100;
    16'b0000000100000010: out_v[220] = 10'b1110110010;
    16'b0010100110000010: out_v[220] = 10'b0100111100;
    16'b0010100100000000: out_v[220] = 10'b1101001101;
    16'b1110101100000000: out_v[220] = 10'b0101101001;
    16'b0010100000000010: out_v[220] = 10'b1101100110;
    16'b1110100100000010: out_v[220] = 10'b1111011011;
    16'b1000100000000010: out_v[220] = 10'b0111011000;
    16'b1010100110000010: out_v[220] = 10'b1101110110;
    16'b0010100000000000: out_v[220] = 10'b1110100010;
    16'b1000100100000010: out_v[220] = 10'b0101011100;
    16'b1100100100000010: out_v[220] = 10'b0100011111;
    16'b0010000000000000: out_v[220] = 10'b0000111000;
    16'b0010000100000000: out_v[220] = 10'b0000110110;
    16'b0010001100000000: out_v[220] = 10'b1101000010;
    16'b0010001000100000: out_v[220] = 10'b0011011000;
    16'b0010000000100000: out_v[220] = 10'b0111011000;
    16'b0000001000100000: out_v[220] = 10'b0011111001;
    16'b0010100000100000: out_v[220] = 10'b1110101010;
    16'b0010001100100000: out_v[220] = 10'b0010111001;
    16'b0010101110100000: out_v[220] = 10'b0010011111;
    16'b1010000100000000: out_v[220] = 10'b0111100101;
    16'b0110100000000010: out_v[220] = 10'b0111100110;
    16'b0010100000100010: out_v[220] = 10'b0010100010;
    16'b1100101000000010: out_v[220] = 10'b1011101101;
    16'b1000101000100010: out_v[220] = 10'b1111001101;
    16'b1010000010000000: out_v[220] = 10'b1111001011;
    16'b1010000000000010: out_v[220] = 10'b0110110111;
    16'b0000101000100010: out_v[220] = 10'b0001101100;
    16'b0000101000000010: out_v[220] = 10'b0001111101;
    16'b0000000000000000: out_v[220] = 10'b1011101010;
    16'b1010000110000000: out_v[220] = 10'b1000110011;
    16'b1000000000000000: out_v[220] = 10'b0010100011;
    16'b1010000000000000: out_v[220] = 10'b1010100111;
    16'b0100101000000010: out_v[220] = 10'b1001010111;
    16'b0000000110000000: out_v[220] = 10'b0001100011;
    16'b0010000110000000: out_v[220] = 10'b0010100011;
    16'b1010001000000000: out_v[220] = 10'b1101001011;
    16'b1000000110000000: out_v[220] = 10'b0011100110;
    16'b1010000000100000: out_v[220] = 10'b1100010110;
    16'b1000001000000000: out_v[220] = 10'b0000110110;
    16'b1000000100000000: out_v[220] = 10'b1011100111;
    16'b1000001000100010: out_v[220] = 10'b0111011011;
    16'b1010001000100010: out_v[220] = 10'b1101001001;
    16'b1010000000100010: out_v[220] = 10'b1001110010;
    16'b0000001100100000: out_v[220] = 10'b0000110111;
    16'b0010000100100000: out_v[220] = 10'b0001001010;
    16'b0000000000100000: out_v[220] = 10'b0001011110;
    16'b1010001000100000: out_v[220] = 10'b1101000010;
    16'b0010000000100010: out_v[220] = 10'b1110110101;
    16'b0000000100100000: out_v[220] = 10'b0101110110;
    16'b0001100000000010: out_v[220] = 10'b0011101110;
    16'b0000100100000010: out_v[220] = 10'b1001010110;
    16'b0011100000000010: out_v[220] = 10'b1010001110;
    16'b0000110000000010: out_v[220] = 10'b1001011011;
    16'b0010110000000010: out_v[220] = 10'b0101010101;
    16'b0010101110000000: out_v[220] = 10'b1100001000;
    16'b1010001100000000: out_v[220] = 10'b0110111010;
    16'b0010101010100010: out_v[220] = 10'b1011100000;
    16'b0010101110100010: out_v[220] = 10'b1011101110;
    default: out_v[220] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000000000110: out_v[221] = 10'b0001100100;
    16'b0000100000000110: out_v[221] = 10'b1010010101;
    16'b0000100001000110: out_v[221] = 10'b1110010001;
    16'b0000100001000010: out_v[221] = 10'b1100100101;
    16'b0000000001000110: out_v[221] = 10'b1011110000;
    16'b0000000000000010: out_v[221] = 10'b0011110100;
    16'b0000000000000100: out_v[221] = 10'b0101011100;
    16'b0000100001000100: out_v[221] = 10'b1111010011;
    16'b0000100001000000: out_v[221] = 10'b1111001110;
    16'b0000100000000010: out_v[221] = 10'b0110100100;
    16'b0000100000000100: out_v[221] = 10'b1000001111;
    16'b0000100000000000: out_v[221] = 10'b0110000010;
    16'b0000000001000010: out_v[221] = 10'b1001111111;
    16'b0000101001000000: out_v[221] = 10'b0100011111;
    16'b0000000000000000: out_v[221] = 10'b1001011111;
    16'b0000101001000110: out_v[221] = 10'b0110111111;
    16'b0100001000000000: out_v[221] = 10'b1000001110;
    16'b0110000000000000: out_v[221] = 10'b1110011101;
    16'b0000001000000000: out_v[221] = 10'b0010011011;
    16'b0110001000000000: out_v[221] = 10'b0101101100;
    16'b0100000000000100: out_v[221] = 10'b1000110101;
    16'b0100000000000000: out_v[221] = 10'b1000111101;
    16'b0100001000000100: out_v[221] = 10'b0000110011;
    16'b0100101000000100: out_v[221] = 10'b0110000100;
    16'b0000001000000010: out_v[221] = 10'b0011001110;
    16'b0000001000000100: out_v[221] = 10'b1011011010;
    16'b0000101000000000: out_v[221] = 10'b1001011110;
    16'b0000100010000000: out_v[221] = 10'b1010100111;
    16'b0110001000000100: out_v[221] = 10'b0110110111;
    16'b0000100010000010: out_v[221] = 10'b0010011100;
    16'b0000101000000100: out_v[221] = 10'b1110011110;
    16'b0000001000000110: out_v[221] = 10'b1010011000;
    16'b0000100010000100: out_v[221] = 10'b1010101011;
    16'b0000101000000110: out_v[221] = 10'b0010001001;
    16'b0100001000000110: out_v[221] = 10'b0100011001;
    16'b0000000010000100: out_v[221] = 10'b1111001101;
    16'b0000000010000000: out_v[221] = 10'b0001001101;
    16'b0000100000001010: out_v[221] = 10'b0100011111;
    16'b0000001001000100: out_v[221] = 10'b0000110010;
    16'b0000000001000000: out_v[221] = 10'b1001110010;
    16'b0000000001000100: out_v[221] = 10'b1100110010;
    16'b0000101001000100: out_v[221] = 10'b1001111001;
    16'b0000001001000000: out_v[221] = 10'b1011110011;
    16'b0000000000001110: out_v[221] = 10'b1110110011;
    16'b0000110000000000: out_v[221] = 10'b0000101000;
    16'b0000110000000010: out_v[221] = 10'b0000100000;
    16'b0000000000001010: out_v[221] = 10'b1011100010;
    16'b0000000000001000: out_v[221] = 10'b0010110000;
    16'b0000000000100110: out_v[221] = 10'b1001100100;
    16'b0000000000100100: out_v[221] = 10'b1001011111;
    16'b0000000000100010: out_v[221] = 10'b0111101100;
    16'b0000000000100000: out_v[221] = 10'b1111001100;
    16'b0000101000000010: out_v[221] = 10'b0110110010;
    default: out_v[221] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0011000010000000: out_v[222] = 10'b1000101100;
    16'b0101000010000000: out_v[222] = 10'b0110110001;
    16'b1010000000000000: out_v[222] = 10'b0001011001;
    16'b0010000000000000: out_v[222] = 10'b1001001100;
    16'b0100000010000000: out_v[222] = 10'b0010110101;
    16'b0110000010000000: out_v[222] = 10'b0010100001;
    16'b0000000010000000: out_v[222] = 10'b1111001111;
    16'b0010000010000000: out_v[222] = 10'b0010011110;
    16'b0100000000000000: out_v[222] = 10'b0011010110;
    16'b0000000010001000: out_v[222] = 10'b1101110001;
    16'b0110000010001000: out_v[222] = 10'b1011101000;
    16'b0100000010001000: out_v[222] = 10'b1001110111;
    16'b1011000000000000: out_v[222] = 10'b0110101011;
    16'b0011000000000000: out_v[222] = 10'b1101001111;
    16'b0111000010000000: out_v[222] = 10'b0110100001;
    16'b1011000010000000: out_v[222] = 10'b0000100001;
    16'b1111000010000000: out_v[222] = 10'b1001100111;
    16'b1000000000000000: out_v[222] = 10'b1010010100;
    16'b0000000000000000: out_v[222] = 10'b0111011011;
    16'b1110000010000000: out_v[222] = 10'b0010100101;
    16'b1010000000100000: out_v[222] = 10'b0111011100;
    16'b0010000000100000: out_v[222] = 10'b1000110011;
    16'b1010000010000000: out_v[222] = 10'b0011110000;
    16'b1001000000000000: out_v[222] = 10'b0100110111;
    16'b0001000010000000: out_v[222] = 10'b0011110100;
    16'b0010000010100000: out_v[222] = 10'b1101001010;
    16'b1110000000000000: out_v[222] = 10'b0001110011;
    16'b0001000000000000: out_v[222] = 10'b0100101111;
    16'b1111000000000000: out_v[222] = 10'b1010110111;
    16'b1000000010000000: out_v[222] = 10'b1000001110;
    16'b0110000000000000: out_v[222] = 10'b0010000111;
    16'b0110000010100000: out_v[222] = 10'b1111110011;
    16'b0001000010001000: out_v[222] = 10'b0100010011;
    16'b0100000000001000: out_v[222] = 10'b0011011000;
    16'b0101000010001000: out_v[222] = 10'b1000000110;
    16'b1000000000001000: out_v[222] = 10'b1110100110;
    16'b0000000000001000: out_v[222] = 10'b0110101110;
    16'b1000000010001000: out_v[222] = 10'b0110011101;
    16'b1100000010001000: out_v[222] = 10'b1100001100;
    16'b1100000000000000: out_v[222] = 10'b1010100010;
    16'b1100000000001000: out_v[222] = 10'b1001101000;
    16'b1110000000001000: out_v[222] = 10'b1101010010;
    16'b1100000010000000: out_v[222] = 10'b1100001110;
    16'b0110000000001000: out_v[222] = 10'b1101011000;
    16'b1110000010001000: out_v[222] = 10'b1010100101;
    16'b1010000010001000: out_v[222] = 10'b1100000010;
    16'b1101000010001000: out_v[222] = 10'b0110011001;
    16'b1101000000001000: out_v[222] = 10'b0001111010;
    16'b1001000010001000: out_v[222] = 10'b1111011000;
    16'b0101000000001000: out_v[222] = 10'b0101001101;
    16'b1001000010000000: out_v[222] = 10'b1010001011;
    16'b1111000010001000: out_v[222] = 10'b1001010110;
    16'b0111000000001000: out_v[222] = 10'b0001011110;
    16'b1111000000001000: out_v[222] = 10'b0101110110;
    16'b1101000010000000: out_v[222] = 10'b1101001111;
    16'b0111000010001000: out_v[222] = 10'b1001001000;
    16'b1011000010001000: out_v[222] = 10'b0001111110;
    16'b0011000000001000: out_v[222] = 10'b0101110111;
    16'b0010000000001000: out_v[222] = 10'b1000101111;
    16'b0111000000000000: out_v[222] = 10'b0110011111;
    16'b0101000000000000: out_v[222] = 10'b0011010100;
    16'b0000000000100000: out_v[222] = 10'b1001010111;
    16'b0100000000100000: out_v[222] = 10'b0111010110;
    16'b1011000000001000: out_v[222] = 10'b0001110011;
    16'b0000000110001000: out_v[222] = 10'b1100111100;
    16'b0011000010001000: out_v[222] = 10'b0111001011;
    16'b1010000000001000: out_v[222] = 10'b1000110010;
    16'b0000000110000000: out_v[222] = 10'b1110001011;
    16'b1001000000001000: out_v[222] = 10'b0001100010;
    16'b0010000010001000: out_v[222] = 10'b0110001001;
    16'b0011000110000000: out_v[222] = 10'b0101010011;
    16'b0001000000001000: out_v[222] = 10'b0100110110;
    16'b0001000110000000: out_v[222] = 10'b1010010110;
    16'b0010000110001000: out_v[222] = 10'b0010101111;
    16'b1101000000000000: out_v[222] = 10'b0011110101;
    16'b0111000010000100: out_v[222] = 10'b1101000100;
    16'b0111000010100000: out_v[222] = 10'b0011001000;
    16'b0110000010000100: out_v[222] = 10'b0111101001;
    16'b0011000010000100: out_v[222] = 10'b0111010001;
    16'b0010000010000100: out_v[222] = 10'b0010101011;
    default: out_v[222] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000110000101000: out_v[223] = 10'b0011001001;
    16'b0000100100111000: out_v[223] = 10'b1010010011;
    16'b0000110100111001: out_v[223] = 10'b0111111011;
    16'b0100110010110001: out_v[223] = 10'b0111011101;
    16'b0000110000100001: out_v[223] = 10'b1110000101;
    16'b0000100100111001: out_v[223] = 10'b1101011101;
    16'b0000110000000001: out_v[223] = 10'b0010100101;
    16'b0100110010010001: out_v[223] = 10'b0111010010;
    16'b0000010000000001: out_v[223] = 10'b1010100010;
    16'b0000110000001000: out_v[223] = 10'b0110100001;
    16'b0100100110111000: out_v[223] = 10'b1101100010;
    16'b0100100110101000: out_v[223] = 10'b0010110111;
    16'b0000110000111001: out_v[223] = 10'b1110001111;
    16'b0000010000101000: out_v[223] = 10'b1110000000;
    16'b0000010000101001: out_v[223] = 10'b1000010101;
    16'b0100110010011001: out_v[223] = 10'b0011110010;
    16'b0100110010111001: out_v[223] = 10'b1101110111;
    16'b0100110110111000: out_v[223] = 10'b1101000001;
    16'b0000110100100001: out_v[223] = 10'b1000110111;
    16'b0100110000101001: out_v[223] = 10'b0010110100;
    16'b0000110000010001: out_v[223] = 10'b1111010010;
    16'b0000000000100001: out_v[223] = 10'b0000111011;
    16'b0000010000111001: out_v[223] = 10'b1101110011;
    16'b0000110000110001: out_v[223] = 10'b0111010111;
    16'b0000100100011000: out_v[223] = 10'b1111100000;
    16'b0000110100110001: out_v[223] = 10'b0010100001;
    16'b0100010010111001: out_v[223] = 10'b1011010011;
    16'b0000110100101000: out_v[223] = 10'b0011010001;
    16'b0100010000101001: out_v[223] = 10'b0100100011;
    16'b0100010010010001: out_v[223] = 10'b0011101101;
    16'b0000010000100001: out_v[223] = 10'b1101000010;
    16'b0000101100111000: out_v[223] = 10'b1011001110;
    16'b0100110010101000: out_v[223] = 10'b1110111111;
    16'b0000010000010001: out_v[223] = 10'b1011011011;
    16'b0000110000101001: out_v[223] = 10'b1000010100;
    16'b0000110100101001: out_v[223] = 10'b1110100111;
    16'b0100110000111001: out_v[223] = 10'b1111001010;
    16'b0000010000110001: out_v[223] = 10'b1001101111;
    16'b0000100100101000: out_v[223] = 10'b1010010011;
    16'b0100010010101001: out_v[223] = 10'b1010011011;
    16'b0000110100001000: out_v[223] = 10'b0110011001;
    16'b0000110100010001: out_v[223] = 10'b1010000111;
    16'b0100110110111001: out_v[223] = 10'b1110001101;
    16'b0100010000100001: out_v[223] = 10'b1000011111;
    16'b0000101100111001: out_v[223] = 10'b1111101111;
    16'b0100111010111001: out_v[223] = 10'b0110011011;
    16'b0000110000011001: out_v[223] = 10'b1111100011;
    16'b0000110000100000: out_v[223] = 10'b0000101011;
    16'b0000010000100000: out_v[223] = 10'b0110000011;
    16'b0100110000101000: out_v[223] = 10'b1000111110;
    16'b0100110010101001: out_v[223] = 10'b1110100111;
    16'b0000110000001001: out_v[223] = 10'b0011111000;
    16'b0000111000111001: out_v[223] = 10'b1000000111;
    16'b0100110110101000: out_v[223] = 10'b0110110110;
    16'b0000000110000000: out_v[223] = 10'b1011000111;
    16'b0000000100000000: out_v[223] = 10'b0101101110;
    16'b0000100100000000: out_v[223] = 10'b0000111100;
    16'b0100000110000000: out_v[223] = 10'b1011101111;
    16'b0000000000000000: out_v[223] = 10'b0100001111;
    16'b0000110100000000: out_v[223] = 10'b1000000110;
    16'b0000000010000000: out_v[223] = 10'b1101001111;
    16'b0100000100000000: out_v[223] = 10'b0010111011;
    16'b0100100110000000: out_v[223] = 10'b0011011010;
    16'b0000000000010000: out_v[223] = 10'b0100010010;
    16'b0000000100010000: out_v[223] = 10'b0011100110;
    16'b0100000010000000: out_v[223] = 10'b0000100111;
    16'b0100000000000000: out_v[223] = 10'b1100100010;
    16'b0100100100000000: out_v[223] = 10'b0111010011;
    16'b0000100000000000: out_v[223] = 10'b1000001001;
    16'b0100000000111000: out_v[223] = 10'b1001110110;
    16'b0000010000000000: out_v[223] = 10'b0011110101;
    16'b0100010100000000: out_v[223] = 10'b0110101101;
    16'b0100000010010000: out_v[223] = 10'b1100000110;
    16'b0100000110010000: out_v[223] = 10'b1011001101;
    16'b0000110000000000: out_v[223] = 10'b0001101001;
    16'b0000000000001000: out_v[223] = 10'b1011100100;
    16'b0100111010111000: out_v[223] = 10'b1001000100;
    16'b0100010010110000: out_v[223] = 10'b1110110011;
    16'b0100011010111000: out_v[223] = 10'b0011001111;
    16'b0100001010111000: out_v[223] = 10'b0001001110;
    16'b0000000000101000: out_v[223] = 10'b0001010110;
    16'b0100010000010000: out_v[223] = 10'b1101011111;
    16'b0000000000111000: out_v[223] = 10'b1010010011;
    16'b0000000000011000: out_v[223] = 10'b1010111110;
    16'b0100010010111000: out_v[223] = 10'b1100100111;
    16'b0000010000111000: out_v[223] = 10'b1011100110;
    16'b0100001010110000: out_v[223] = 10'b0111110101;
    16'b0100000000010000: out_v[223] = 10'b1110110101;
    16'b0100010000000000: out_v[223] = 10'b1001110011;
    16'b0000010000011000: out_v[223] = 10'b0001111110;
    16'b0100010010000000: out_v[223] = 10'b0010111010;
    16'b0100010010010000: out_v[223] = 10'b1100010110;
    16'b0100000000101000: out_v[223] = 10'b1101110010;
    16'b0000010000001000: out_v[223] = 10'b0011001011;
    16'b0100000010110000: out_v[223] = 10'b0110110111;
    16'b0000111000111000: out_v[223] = 10'b0001011110;
    16'b0000010100000000: out_v[223] = 10'b1101000000;
    16'b0100000010111000: out_v[223] = 10'b0011110111;
    16'b0000010000010000: out_v[223] = 10'b1001101101;
    16'b0100001010010000: out_v[223] = 10'b1110000010;
    16'b0100011010110000: out_v[223] = 10'b1110111101;
    16'b0100110010111000: out_v[223] = 10'b1000111110;
    16'b0100110010010000: out_v[223] = 10'b1011110011;
    16'b0100000010101000: out_v[223] = 10'b1100100111;
    16'b0000110000111000: out_v[223] = 10'b1111001110;
    16'b0000010100011000: out_v[223] = 10'b0111000011;
    16'b0100000110011000: out_v[223] = 10'b1010010111;
    16'b0000100100001000: out_v[223] = 10'b0000111001;
    16'b0100001110111000: out_v[223] = 10'b0110011111;
    16'b0000000100001000: out_v[223] = 10'b0111100001;
    16'b0100000100011000: out_v[223] = 10'b0111101000;
    16'b0000010100001000: out_v[223] = 10'b0001101001;
    16'b0100011110011000: out_v[223] = 10'b1111011111;
    16'b0000000100011000: out_v[223] = 10'b1111010000;
    16'b0000110100111000: out_v[223] = 10'b1111011110;
    16'b0000011100111000: out_v[223] = 10'b1110011010;
    16'b0000110100011000: out_v[223] = 10'b0101001100;
    16'b0000001100011000: out_v[223] = 10'b1111011001;
    16'b0100001110011000: out_v[223] = 10'b1010001101;
    16'b0000110100001001: out_v[223] = 10'b1110101000;
    16'b0100010110011000: out_v[223] = 10'b1010001011;
    16'b0000011100011000: out_v[223] = 10'b0111001011;
    16'b0000100100001001: out_v[223] = 10'b0110011100;
    16'b0000000100001001: out_v[223] = 10'b1111100111;
    16'b0100001110010000: out_v[223] = 10'b0001011001;
    16'b0000010100010000: out_v[223] = 10'b0101001001;
    16'b0000010100111000: out_v[223] = 10'b0111110110;
    16'b0100000100001000: out_v[223] = 10'b1110111001;
    16'b0000110100100000: out_v[223] = 10'b0111001001;
    16'b0000111100111000: out_v[223] = 10'b1001110010;
    16'b0000000000001001: out_v[223] = 10'b0000110010;
    16'b0000010000001001: out_v[223] = 10'b0100011001;
    16'b0100000010001001: out_v[223] = 10'b1111001011;
    16'b0000010100001001: out_v[223] = 10'b1100110110;
    16'b0000000000000001: out_v[223] = 10'b0000110001;
    16'b0000000100101001: out_v[223] = 10'b0111000100;
    16'b0000000000101001: out_v[223] = 10'b0101011001;
    16'b0000100000101000: out_v[223] = 10'b1100001011;
    16'b0000100100100000: out_v[223] = 10'b1110110000;
    16'b0000100000001000: out_v[223] = 10'b0110001011;
    16'b0000010100101001: out_v[223] = 10'b1101010110;
    16'b0000100000001001: out_v[223] = 10'b0101001011;
    16'b0000000100000001: out_v[223] = 10'b1011100000;
    16'b0000100000101001: out_v[223] = 10'b1100010110;
    16'b0000010100000001: out_v[223] = 10'b1101100010;
    16'b0000000100110000: out_v[223] = 10'b1001100111;
    16'b0000100100010000: out_v[223] = 10'b0111010001;
    16'b0000110100011001: out_v[223] = 10'b0001100111;
    16'b0000110100000001: out_v[223] = 10'b1111000000;
    16'b0000100000010000: out_v[223] = 10'b0101011001;
    16'b0000110100010000: out_v[223] = 10'b1111110011;
    16'b0000110000010000: out_v[223] = 10'b0101011001;
    16'b0000100000000001: out_v[223] = 10'b0111110100;
    16'b0000000100100000: out_v[223] = 10'b0111100000;
    16'b0000010100011001: out_v[223] = 10'b0111100000;
    16'b0000100100000001: out_v[223] = 10'b0110011110;
    16'b0100010110001001: out_v[223] = 10'b1011100011;
    16'b0100010110001000: out_v[223] = 10'b0010111101;
    16'b0100010110011001: out_v[223] = 10'b1110110111;
    16'b0100110110011000: out_v[223] = 10'b1110110111;
    16'b0100110110001000: out_v[223] = 10'b1100100100;
    16'b0100110010001000: out_v[223] = 10'b1001001111;
    16'b0100110100001000: out_v[223] = 10'b1111100000;
    16'b0100110110001001: out_v[223] = 10'b1011011010;
    16'b0100100110001000: out_v[223] = 10'b1101001010;
    16'b0000100110001000: out_v[223] = 10'b1011010010;
    16'b0100110110000000: out_v[223] = 10'b1100011001;
    16'b0100010010001001: out_v[223] = 10'b1011001011;
    16'b0100110000001001: out_v[223] = 10'b1111100000;
    16'b0100100010001000: out_v[223] = 10'b0011101001;
    16'b0100100100001000: out_v[223] = 10'b1101010111;
    16'b0100100010000000: out_v[223] = 10'b0000011101;
    16'b0100010000001001: out_v[223] = 10'b1111011011;
    16'b0000000000100000: out_v[223] = 10'b1001101111;
    16'b0100100000001000: out_v[223] = 10'b0111001011;
    16'b0000010100100001: out_v[223] = 10'b0111100000;
    16'b0100110010001001: out_v[223] = 10'b0101111011;
    16'b0100110010000000: out_v[223] = 10'b1001100100;
    16'b0000000100100001: out_v[223] = 10'b0111100011;
    16'b0100110000001000: out_v[223] = 10'b0010101111;
    16'b0100010000001000: out_v[223] = 10'b1011011011;
    16'b0100100110011000: out_v[223] = 10'b1110110001;
    16'b0000100100101001: out_v[223] = 10'b0100111110;
    16'b0000100000100001: out_v[223] = 10'b0111100010;
    16'b0000110000101010: out_v[223] = 10'b0111011010;
    16'b0000110000000010: out_v[223] = 10'b0011100111;
    16'b0000110000001011: out_v[223] = 10'b1111011010;
    16'b0000100000100000: out_v[223] = 10'b1101000110;
    16'b0000110000101011: out_v[223] = 10'b0110100110;
    16'b0000110000001010: out_v[223] = 10'b1111000111;
    16'b0000110100110000: out_v[223] = 10'b0101100111;
    16'b0000010100110000: out_v[223] = 10'b1110100101;
    16'b0100110110100000: out_v[223] = 10'b1100111011;
    16'b0100100110100000: out_v[223] = 10'b1111001010;
    16'b0000100100110000: out_v[223] = 10'b0101000101;
    16'b0000110000110000: out_v[223] = 10'b0011111111;
    16'b0100010110000000: out_v[223] = 10'b1100100001;
    16'b0000010100100000: out_v[223] = 10'b0001110111;
    16'b0100110100000000: out_v[223] = 10'b0011001101;
    16'b0000010100101000: out_v[223] = 10'b1001010010;
    16'b0000110100000011: out_v[223] = 10'b1000101011;
    16'b0000110000000011: out_v[223] = 10'b1000101010;
    16'b0000010000000011: out_v[223] = 10'b1011100111;
    default: out_v[223] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000010100010011: out_v[224] = 10'b1001101101;
    16'b0100110000000011: out_v[224] = 10'b0101110010;
    16'b0000110000010011: out_v[224] = 10'b0101000101;
    16'b0000110000000000: out_v[224] = 10'b0110010110;
    16'b0100110000000000: out_v[224] = 10'b1110000011;
    16'b0100110000010011: out_v[224] = 10'b0110001001;
    16'b0100110000010010: out_v[224] = 10'b0011001111;
    16'b0000110100000011: out_v[224] = 10'b1001101101;
    16'b0000110000000011: out_v[224] = 10'b0111011011;
    16'b0000110100010011: out_v[224] = 10'b1001001010;
    16'b0000110010010011: out_v[224] = 10'b0110000011;
    16'b0000110000010000: out_v[224] = 10'b0111010001;
    16'b0000100000000000: out_v[224] = 10'b0111010000;
    16'b0000110001010011: out_v[224] = 10'b1100100001;
    16'b0000010000000011: out_v[224] = 10'b1000111011;
    16'b0000110101010011: out_v[224] = 10'b0111111011;
    16'b0100110100000000: out_v[224] = 10'b1010001110;
    16'b0000010100010000: out_v[224] = 10'b1110010100;
    16'b0000110011010011: out_v[224] = 10'b0011011100;
    16'b0000010100000011: out_v[224] = 10'b0011001000;
    16'b0100100000000000: out_v[224] = 10'b1111011111;
    16'b0000010100000000: out_v[224] = 10'b1101000011;
    16'b0100110100010011: out_v[224] = 10'b1101100111;
    16'b0000000100010011: out_v[224] = 10'b0100101001;
    16'b0000010000010011: out_v[224] = 10'b0000001110;
    16'b0100110001010011: out_v[224] = 10'b1111001010;
    16'b0000100000010011: out_v[224] = 10'b0101010101;
    16'b0000100000010000: out_v[224] = 10'b0111100111;
    16'b0100110000000010: out_v[224] = 10'b1111110111;
    16'b0000010100010001: out_v[224] = 10'b1110010101;
    16'b0000000100000000: out_v[224] = 10'b1011101111;
    16'b0100110100000011: out_v[224] = 10'b1010000011;
    16'b0000110110010011: out_v[224] = 10'b0011000101;
    16'b0000100001010000: out_v[224] = 10'b0101001101;
    16'b0000010001010011: out_v[224] = 10'b1010111000;
    16'b0100110000010000: out_v[224] = 10'b0000001011;
    16'b0000000000000000: out_v[224] = 10'b1000101010;
    16'b0000010000010000: out_v[224] = 10'b1101100011;
    16'b0000000000010000: out_v[224] = 10'b1010011000;
    16'b0000010000000001: out_v[224] = 10'b0110111001;
    16'b0000010000010001: out_v[224] = 10'b1000001111;
    16'b0000010000000000: out_v[224] = 10'b1101110000;
    16'b0000010010010001: out_v[224] = 10'b0111011001;
    16'b0000010010010011: out_v[224] = 10'b1001101011;
    16'b0100000100000000: out_v[224] = 10'b0110011010;
    16'b0000010110010011: out_v[224] = 10'b1100110100;
    16'b0000010101010011: out_v[224] = 10'b0000111110;
    16'b0000000100010000: out_v[224] = 10'b0110010100;
    16'b0000000100010010: out_v[224] = 10'b1110110110;
    16'b0000010110010000: out_v[224] = 10'b1110111011;
    16'b0000100100000000: out_v[224] = 10'b1001101101;
    16'b0000010110010001: out_v[224] = 10'b1011110110;
    16'b0000000110000000: out_v[224] = 10'b1011001001;
    16'b0100000100010000: out_v[224] = 10'b0110100010;
    16'b0000010111010011: out_v[224] = 10'b1011101000;
    16'b0000000110010000: out_v[224] = 10'b1000110111;
    16'b0000000110010010: out_v[224] = 10'b1111011100;
    16'b0000000101000000: out_v[224] = 10'b0000100110;
    16'b0000000101010000: out_v[224] = 10'b1100010111;
    16'b0000000101010010: out_v[224] = 10'b1101011110;
    16'b0000100100010000: out_v[224] = 10'b1001000111;
    16'b0100000100010011: out_v[224] = 10'b1011010011;
    16'b0000000100000010: out_v[224] = 10'b1011010101;
    16'b0000010110010010: out_v[224] = 10'b1011100101;
    16'b0100010100010011: out_v[224] = 10'b1101010100;
    16'b0000010110000011: out_v[224] = 10'b1011101010;
    16'b0000010010000011: out_v[224] = 10'b0001111010;
    16'b0000100101010000: out_v[224] = 10'b1111001000;
    16'b0000010100010010: out_v[224] = 10'b1000110110;
    16'b0000100100010011: out_v[224] = 10'b1000110010;
    16'b0000000100000011: out_v[224] = 10'b0010111110;
    16'b0100000100010010: out_v[224] = 10'b0110101111;
    16'b0000000110010011: out_v[224] = 10'b1111010110;
    16'b0000000110000010: out_v[224] = 10'b1111100111;
    16'b0000000111010000: out_v[224] = 10'b0011111010;
    16'b0100010000010000: out_v[224] = 10'b0000111110;
    16'b0000000000010011: out_v[224] = 10'b1001001000;
    16'b0000010010010000: out_v[224] = 10'b0000001101;
    16'b0000000000000011: out_v[224] = 10'b1001011110;
    16'b0100010000010011: out_v[224] = 10'b1001101100;
    16'b0000000000010010: out_v[224] = 10'b1111100010;
    16'b0100000000000000: out_v[224] = 10'b1011111000;
    16'b0100010000000000: out_v[224] = 10'b0000110000;
    16'b0000000000010001: out_v[224] = 10'b0100011100;
    16'b0000100000000011: out_v[224] = 10'b0110110100;
    16'b0000100100000011: out_v[224] = 10'b1000011000;
    16'b0100100100010000: out_v[224] = 10'b1010110011;
    16'b0000010100000001: out_v[224] = 10'b0111010010;
    16'b0100110100000001: out_v[224] = 10'b0111111111;
    16'b0100100100000000: out_v[224] = 10'b1000111001;
    16'b0000110100000000: out_v[224] = 10'b1101110010;
    16'b0000100100000010: out_v[224] = 10'b0000011010;
    16'b0000110000000001: out_v[224] = 10'b0101011110;
    16'b0000110100010000: out_v[224] = 10'b1001110110;
    16'b0100100000010000: out_v[224] = 10'b0110110111;
    16'b0000110100010001: out_v[224] = 10'b0111110010;
    16'b0100110100010000: out_v[224] = 10'b0100011001;
    16'b0000110100000001: out_v[224] = 10'b1000000101;
    16'b0000100000000010: out_v[224] = 10'b0100110111;
    16'b0100100100000011: out_v[224] = 10'b0001110110;
    16'b0100010000000011: out_v[224] = 10'b1001001010;
    16'b0100010100000000: out_v[224] = 10'b0110000111;
    16'b0100010100000011: out_v[224] = 10'b1101001101;
    16'b0100010000000001: out_v[224] = 10'b0111000101;
    16'b0100010000010001: out_v[224] = 10'b0001101110;
    16'b0100000000010011: out_v[224] = 10'b1111100110;
    16'b0000110101000011: out_v[224] = 10'b0111001011;
    16'b0000110111000011: out_v[224] = 10'b0101010010;
    16'b0000110100010010: out_v[224] = 10'b0111101100;
    16'b0000110111010011: out_v[224] = 10'b1101110110;
    16'b0000010100000010: out_v[224] = 10'b1001111011;
    16'b0000110010000011: out_v[224] = 10'b0011110111;
    16'b1000010100000000: out_v[224] = 10'b1110011111;
    16'b0000100100010010: out_v[224] = 10'b1001000011;
    16'b1000010100000011: out_v[224] = 10'b1010110011;
    16'b1000000100000000: out_v[224] = 10'b0101111010;
    16'b0000110110000011: out_v[224] = 10'b1010011001;
    16'b0000010000000100: out_v[224] = 10'b0111010101;
    16'b0000000000000100: out_v[224] = 10'b1010011110;
    16'b0100010100010001: out_v[224] = 10'b1011100111;
    16'b0100010100010000: out_v[224] = 10'b1100000011;
    16'b0100010100000001: out_v[224] = 10'b0001111111;
    default: out_v[224] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1010100000000000: out_v[225] = 10'b1000111001;
    16'b0010100010001000: out_v[225] = 10'b1100001111;
    16'b1010100010001000: out_v[225] = 10'b1100001001;
    16'b1000000010001000: out_v[225] = 10'b1000110001;
    16'b0010000010001000: out_v[225] = 10'b0110001101;
    16'b1010000000000000: out_v[225] = 10'b0111100110;
    16'b1010100010000000: out_v[225] = 10'b1001100101;
    16'b0010100000000000: out_v[225] = 10'b1010000010;
    16'b1010100000001000: out_v[225] = 10'b1110000010;
    16'b0000100010001000: out_v[225] = 10'b1110001011;
    16'b1010000010001000: out_v[225] = 10'b0110001001;
    16'b1010100010001001: out_v[225] = 10'b0011111011;
    16'b0010100010000000: out_v[225] = 10'b1100110001;
    16'b1010000010001001: out_v[225] = 10'b1010011111;
    16'b1010000010000000: out_v[225] = 10'b0010110110;
    16'b0000000010001000: out_v[225] = 10'b0000111011;
    16'b0010000000001000: out_v[225] = 10'b1000010011;
    16'b0010000000000000: out_v[225] = 10'b0111011001;
    16'b1000000000000000: out_v[225] = 10'b0101000011;
    16'b0010100000001000: out_v[225] = 10'b1011001000;
    16'b0010000010000000: out_v[225] = 10'b0110011000;
    16'b1000100000000000: out_v[225] = 10'b0011011110;
    16'b1010100000000101: out_v[225] = 10'b0010111011;
    16'b1010100000000001: out_v[225] = 10'b1111001001;
    16'b1010100010000001: out_v[225] = 10'b1110000111;
    16'b1000100010001000: out_v[225] = 10'b1101001011;
    16'b1010000000001000: out_v[225] = 10'b0101000001;
    16'b0000000000000000: out_v[225] = 10'b1000001111;
    16'b0000000000000001: out_v[225] = 10'b1001011010;
    16'b1000000000000001: out_v[225] = 10'b0100101111;
    16'b1000000000100101: out_v[225] = 10'b0110011101;
    16'b1010100010000101: out_v[225] = 10'b1011011010;
    16'b1000000000000101: out_v[225] = 10'b1101111100;
    16'b1010000000100101: out_v[225] = 10'b1100101011;
    16'b1010000000000101: out_v[225] = 10'b0010111010;
    16'b1000100010000000: out_v[225] = 10'b1001000100;
    16'b1010000010000001: out_v[225] = 10'b0011011111;
    16'b1010000010100101: out_v[225] = 10'b1110000000;
    16'b1000000000100100: out_v[225] = 10'b0101111100;
    16'b1010100010101101: out_v[225] = 10'b1100000111;
    16'b1010000000000001: out_v[225] = 10'b1000110100;
    16'b1010100010100101: out_v[225] = 10'b0111000100;
    16'b1110100010001000: out_v[225] = 10'b1010111111;
    16'b1000000010000000: out_v[225] = 10'b1100110110;
    16'b1010000010010000: out_v[225] = 10'b1010100111;
    16'b1000000000010000: out_v[225] = 10'b1010001100;
    16'b1010000000000100: out_v[225] = 10'b1110110111;
    16'b1010100000100101: out_v[225] = 10'b1100100101;
    16'b1010000010000101: out_v[225] = 10'b1111100001;
    16'b0000000010000000: out_v[225] = 10'b0101100010;
    16'b1000000000110101: out_v[225] = 10'b0001001001;
    16'b1010000000100100: out_v[225] = 10'b1100110010;
    16'b0000000000100101: out_v[225] = 10'b1101100101;
    16'b0000000000100100: out_v[225] = 10'b0011000111;
    16'b0010000000100100: out_v[225] = 10'b1101111000;
    16'b0010000010100101: out_v[225] = 10'b1111111110;
    16'b1000100000100100: out_v[225] = 10'b1011100101;
    16'b0010000000100101: out_v[225] = 10'b1011001011;
    16'b1110000010000000: out_v[225] = 10'b1011011011;
    16'b0010100000100100: out_v[225] = 10'b0101100001;
    16'b0000000000000100: out_v[225] = 10'b0100111001;
    16'b0010000010100100: out_v[225] = 10'b0100110011;
    16'b1110100010000000: out_v[225] = 10'b0111110011;
    16'b0110000000000000: out_v[225] = 10'b0011011001;
    16'b0000000000000101: out_v[225] = 10'b1101110100;
    16'b0010000000000100: out_v[225] = 10'b1000111010;
    16'b0010000000000001: out_v[225] = 10'b0110111001;
    16'b0010000000000101: out_v[225] = 10'b1101001011;
    16'b0010000010000001: out_v[225] = 10'b0110110101;
    16'b0010100010100100: out_v[225] = 10'b0011111011;
    16'b1000100000100101: out_v[225] = 10'b1110011000;
    16'b0000100000001000: out_v[225] = 10'b0110011010;
    16'b1000100000001000: out_v[225] = 10'b0010011000;
    16'b0000100000000000: out_v[225] = 10'b1110001000;
    16'b0000100000100100: out_v[225] = 10'b0000110111;
    16'b1000000000001000: out_v[225] = 10'b0111101111;
    16'b0000100000101100: out_v[225] = 10'b0010010000;
    16'b0000100010000000: out_v[225] = 10'b0010110111;
    16'b0010100000000100: out_v[225] = 10'b1110100010;
    16'b0000000000001000: out_v[225] = 10'b0001100000;
    16'b1000000000000010: out_v[225] = 10'b1010101001;
    16'b1000100000000010: out_v[225] = 10'b1010001110;
    16'b1000100000000001: out_v[225] = 10'b0011100011;
    16'b1010000000000010: out_v[225] = 10'b0111011010;
    16'b1000100100000001: out_v[225] = 10'b1101000010;
    16'b1000100010000010: out_v[225] = 10'b1111010010;
    16'b1000000000101100: out_v[225] = 10'b1011000010;
    16'b1010100010000010: out_v[225] = 10'b1011001110;
    16'b1000100000000101: out_v[225] = 10'b0011000111;
    16'b1000100010000001: out_v[225] = 10'b0101011010;
    16'b1010000010000010: out_v[225] = 10'b1101010011;
    16'b1000100100000101: out_v[225] = 10'b1111110101;
    default: out_v[225] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1100101100000010: out_v[226] = 10'b1011001111;
    16'b1000100100000010: out_v[226] = 10'b1001001101;
    16'b1000101100000010: out_v[226] = 10'b1010011111;
    16'b1000000100000000: out_v[226] = 10'b1010001101;
    16'b1000000110000010: out_v[226] = 10'b1111001100;
    16'b1000100100000000: out_v[226] = 10'b1010000000;
    16'b1000000000000000: out_v[226] = 10'b0010100011;
    16'b0000001000000010: out_v[226] = 10'b1000111011;
    16'b0000001010000010: out_v[226] = 10'b0011100111;
    16'b1000000000000010: out_v[226] = 10'b0101011010;
    16'b0000100100000010: out_v[226] = 10'b0111110100;
    16'b0000100100000000: out_v[226] = 10'b1011000100;
    16'b0000101100000010: out_v[226] = 10'b0001101000;
    16'b1000000100000010: out_v[226] = 10'b1111101010;
    16'b1100100100000010: out_v[226] = 10'b0011111100;
    16'b1000101110000010: out_v[226] = 10'b0110010111;
    16'b0000101100000000: out_v[226] = 10'b1001110100;
    16'b1000001110000010: out_v[226] = 10'b1110000101;
    16'b1000001100000010: out_v[226] = 10'b1100001000;
    16'b1000000010000010: out_v[226] = 10'b0111001001;
    16'b1100001010000010: out_v[226] = 10'b0110111011;
    16'b1000001010000010: out_v[226] = 10'b0110011110;
    16'b1000001000000010: out_v[226] = 10'b0101010000;
    16'b0000000100000000: out_v[226] = 10'b1011010110;
    16'b0000001100000010: out_v[226] = 10'b1101000001;
    16'b1000100110000010: out_v[226] = 10'b0100001111;
    16'b0000000000000000: out_v[226] = 10'b1101110001;
    16'b0000000000000010: out_v[226] = 10'b1110100010;
    16'b1000000010000000: out_v[226] = 10'b1001000100;
    16'b0000000010000010: out_v[226] = 10'b1100100111;
    16'b1100001100000010: out_v[226] = 10'b1011000010;
    16'b0000000100000010: out_v[226] = 10'b1100100010;
    16'b1000101100000000: out_v[226] = 10'b1000101001;
    16'b0100000000000010: out_v[226] = 10'b1001010111;
    16'b0000001000000000: out_v[226] = 10'b1010011110;
    16'b0100001000000010: out_v[226] = 10'b1011001110;
    16'b1000101110000000: out_v[226] = 10'b1000010110;
    16'b1000001000000000: out_v[226] = 10'b0011011110;
    16'b0000000010000000: out_v[226] = 10'b0100000111;
    16'b0000001010000000: out_v[226] = 10'b0001000110;
    16'b0000001100000000: out_v[226] = 10'b1001001110;
    16'b1000001010000000: out_v[226] = 10'b1010001001;
    16'b1000001110000000: out_v[226] = 10'b1111111100;
    16'b0000101110000000: out_v[226] = 10'b1101000000;
    16'b1000001100000000: out_v[226] = 10'b0111010110;
    16'b1100001000000010: out_v[226] = 10'b1011101110;
    16'b1000100110000000: out_v[226] = 10'b0100111111;
    16'b0100001100000010: out_v[226] = 10'b1010100101;
    16'b1100000000000010: out_v[226] = 10'b0011111101;
    16'b0100000000000000: out_v[226] = 10'b0100101011;
    16'b0000101110000010: out_v[226] = 10'b0101110000;
    16'b0100101100000010: out_v[226] = 10'b0110111000;
    16'b0101000000000010: out_v[226] = 10'b1000111101;
    16'b0100100100000010: out_v[226] = 10'b1010110110;
    16'b1100000100000010: out_v[226] = 10'b1000101000;
    16'b1001100100000000: out_v[226] = 10'b0011111111;
    16'b0100000100000010: out_v[226] = 10'b0111111110;
    16'b0010000000000000: out_v[226] = 10'b0100111100;
    16'b1010000000000000: out_v[226] = 10'b1101101000;
    16'b1010000000000010: out_v[226] = 10'b1010110010;
    16'b0110000000000010: out_v[226] = 10'b0110011010;
    16'b0100101110000010: out_v[226] = 10'b0011110110;
    16'b1110000000000010: out_v[226] = 10'b1000110111;
    16'b0010000000000010: out_v[226] = 10'b1000111011;
    16'b0000100110000010: out_v[226] = 10'b0111101011;
    16'b0000100110000000: out_v[226] = 10'b1001101011;
    16'b0000001110000000: out_v[226] = 10'b1011010010;
    16'b0000000110000000: out_v[226] = 10'b1010011011;
    16'b0101100100000010: out_v[226] = 10'b0111000010;
    16'b1101000000000010: out_v[226] = 10'b0010011000;
    16'b1101000100000010: out_v[226] = 10'b1111001011;
    16'b1101100100000010: out_v[226] = 10'b0011010110;
    16'b1001100100000010: out_v[226] = 10'b1101110111;
    16'b1001000000000000: out_v[226] = 10'b1101101010;
    16'b1001000000000010: out_v[226] = 10'b0010101010;
    16'b1100000000000000: out_v[226] = 10'b1101010111;
    16'b0100001000000000: out_v[226] = 10'b0101100001;
    16'b1100001000000000: out_v[226] = 10'b0101111100;
    default: out_v[226] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100000001000010: out_v[227] = 10'b1111000011;
    16'b0010000001001010: out_v[227] = 10'b0011011011;
    16'b0110000001001010: out_v[227] = 10'b1011100010;
    16'b0000000001000010: out_v[227] = 10'b1000100011;
    16'b1010000000001010: out_v[227] = 10'b1111110110;
    16'b1010000001001000: out_v[227] = 10'b0011101101;
    16'b1010000000000000: out_v[227] = 10'b1101011011;
    16'b0010000101001010: out_v[227] = 10'b0111000101;
    16'b0000000101001010: out_v[227] = 10'b0001111100;
    16'b0100000001001010: out_v[227] = 10'b1100001111;
    16'b0010000000001010: out_v[227] = 10'b1001000011;
    16'b0000000001001010: out_v[227] = 10'b1010110010;
    16'b1110000001001010: out_v[227] = 10'b0111011110;
    16'b1010000000000010: out_v[227] = 10'b1111011011;
    16'b1100000001001010: out_v[227] = 10'b0110001101;
    16'b1110000001001110: out_v[227] = 10'b1000100001;
    16'b0000000101000010: out_v[227] = 10'b0010011100;
    16'b0010000000000010: out_v[227] = 10'b0011101011;
    16'b1110000000000110: out_v[227] = 10'b0110100011;
    16'b1110000000001010: out_v[227] = 10'b0111111111;
    16'b1010000001001010: out_v[227] = 10'b0101000010;
    16'b1100000001001110: out_v[227] = 10'b1011010011;
    16'b0000000100000010: out_v[227] = 10'b1100111001;
    16'b0010000001001000: out_v[227] = 10'b0100101111;
    16'b0000000000000010: out_v[227] = 10'b0110101111;
    16'b1110000000000010: out_v[227] = 10'b1111110110;
    16'b0010000000000000: out_v[227] = 10'b1000110110;
    16'b0100000001001110: out_v[227] = 10'b0001001100;
    16'b1000000001001000: out_v[227] = 10'b0110111001;
    16'b0100000000000010: out_v[227] = 10'b0001110110;
    16'b0010000101001000: out_v[227] = 10'b0010000101;
    16'b1010000101001010: out_v[227] = 10'b1100110011;
    16'b0110000000000010: out_v[227] = 10'b1100110000;
    16'b0000000100000000: out_v[227] = 10'b1001110001;
    16'b0000000000000000: out_v[227] = 10'b1010000110;
    16'b0100000100000000: out_v[227] = 10'b0100000000;
    16'b0100000100000001: out_v[227] = 10'b1011001110;
    16'b0100001010000111: out_v[227] = 10'b1110001000;
    16'b0000000000000011: out_v[227] = 10'b0100011110;
    16'b0100000100000110: out_v[227] = 10'b1010001111;
    16'b0000000001000000: out_v[227] = 10'b0001110110;
    16'b0010000001000010: out_v[227] = 10'b0001110111;
    16'b0000000001000011: out_v[227] = 10'b1111100100;
    16'b0100000010000110: out_v[227] = 10'b0000111111;
    16'b0100000000000100: out_v[227] = 10'b0111101000;
    16'b0000001010000011: out_v[227] = 10'b1111111011;
    16'b0110000001001100: out_v[227] = 10'b1011011010;
    16'b0110000001001000: out_v[227] = 10'b0010011101;
    16'b0000000101000000: out_v[227] = 10'b1010101111;
    16'b0010000001001001: out_v[227] = 10'b1110110001;
    16'b0100001110000111: out_v[227] = 10'b0001001001;
    16'b0100000010000111: out_v[227] = 10'b1111100011;
    16'b0100000000000110: out_v[227] = 10'b0001011110;
    16'b0010000001000000: out_v[227] = 10'b0111010110;
    16'b0000000101001000: out_v[227] = 10'b1010100110;
    16'b0100000100000010: out_v[227] = 10'b1011100011;
    16'b0010000001001100: out_v[227] = 10'b1011011011;
    16'b0000001000000011: out_v[227] = 10'b1110110101;
    16'b0000000100000011: out_v[227] = 10'b1110011001;
    16'b0000000010000011: out_v[227] = 10'b1001101101;
    16'b0010000101000000: out_v[227] = 10'b1111000011;
    16'b0000000001001000: out_v[227] = 10'b1001011000;
    16'b0110000001000100: out_v[227] = 10'b0110101011;
    16'b0100001010000110: out_v[227] = 10'b0001110110;
    16'b0100001110000110: out_v[227] = 10'b0010111001;
    16'b0010000100000010: out_v[227] = 10'b1001111000;
    16'b0110000100000010: out_v[227] = 10'b0110011000;
    16'b0000001110000011: out_v[227] = 10'b1111110101;
    16'b0100001110000010: out_v[227] = 10'b1101001111;
    16'b0100000110000010: out_v[227] = 10'b1110011011;
    16'b0100001110000000: out_v[227] = 10'b1100011101;
    16'b0100000100000100: out_v[227] = 10'b0100010011;
    16'b0100000110000000: out_v[227] = 10'b1011001011;
    16'b0100000110000110: out_v[227] = 10'b0001011100;
    16'b0000000110000010: out_v[227] = 10'b0001011100;
    16'b0000001110000010: out_v[227] = 10'b1101101111;
    16'b0100001110000100: out_v[227] = 10'b0100011010;
    16'b0000000110000000: out_v[227] = 10'b0001011011;
    16'b0100001100000011: out_v[227] = 10'b1011000001;
    16'b0110001110000011: out_v[227] = 10'b1111101011;
    16'b0100001110000011: out_v[227] = 10'b1110001011;
    16'b0100000100000011: out_v[227] = 10'b0010110001;
    16'b0010000100000011: out_v[227] = 10'b1011111011;
    16'b0100000000000000: out_v[227] = 10'b1110011001;
    16'b0100000101000010: out_v[227] = 10'b0111010010;
    16'b0010000100000000: out_v[227] = 10'b0110101010;
    16'b0100000110000100: out_v[227] = 10'b1101000001;
    16'b0100000110000011: out_v[227] = 10'b0111000000;
    16'b0100000001000000: out_v[227] = 10'b1010111000;
    16'b0100001011001100: out_v[227] = 10'b0100000111;
    16'b0100000001001000: out_v[227] = 10'b1110010010;
    16'b0100000101000000: out_v[227] = 10'b1001011000;
    16'b1000000001001010: out_v[227] = 10'b1011111010;
    16'b0100000101001000: out_v[227] = 10'b1000001111;
    16'b0100000101001100: out_v[227] = 10'b1110011111;
    16'b0100000001000100: out_v[227] = 10'b1001111001;
    16'b0000000001001100: out_v[227] = 10'b1111011010;
    16'b0100000001001100: out_v[227] = 10'b0001011000;
    16'b0100000101000110: out_v[227] = 10'b0111100110;
    16'b0010000101000010: out_v[227] = 10'b0100110001;
    16'b0100000101001010: out_v[227] = 10'b0101010110;
    16'b1000000001000001: out_v[227] = 10'b1110101111;
    16'b1000000001000000: out_v[227] = 10'b0010010011;
    16'b0000000000000001: out_v[227] = 10'b1101100010;
    16'b1000000001001001: out_v[227] = 10'b1110011101;
    16'b1000000101001000: out_v[227] = 10'b0101111111;
    16'b0000010101000000: out_v[227] = 10'b0110111000;
    16'b0000000001000001: out_v[227] = 10'b0001101001;
    16'b0000000001001001: out_v[227] = 10'b1100101110;
    16'b0000010001000000: out_v[227] = 10'b0010110011;
    16'b0000000010000000: out_v[227] = 10'b0110000001;
    16'b0000000010000010: out_v[227] = 10'b0100010110;
    default: out_v[227] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000100011100: out_v[228] = 10'b1100110000;
    16'b0000000000011000: out_v[228] = 10'b1001111100;
    16'b0000001000011000: out_v[228] = 10'b1010001110;
    16'b0000000100011000: out_v[228] = 10'b1101110110;
    16'b0000010000011100: out_v[228] = 10'b0110011110;
    16'b0000001000010000: out_v[228] = 10'b1001000101;
    16'b0000010000011000: out_v[228] = 10'b0110001011;
    16'b0000011000010000: out_v[228] = 10'b1001101011;
    16'b0000000000001100: out_v[228] = 10'b0010010111;
    16'b0000000000001000: out_v[228] = 10'b0000011111;
    16'b0000010100011100: out_v[228] = 10'b1101010011;
    16'b0000000000011100: out_v[228] = 10'b0010111101;
    16'b0000001000110000: out_v[228] = 10'b1110001011;
    16'b0000001000011100: out_v[228] = 10'b1101100000;
    16'b0000011000011000: out_v[228] = 10'b1010001101;
    16'b0000000000111000: out_v[228] = 10'b0010011110;
    16'b0000001000100000: out_v[228] = 10'b1101111001;
    16'b0010001000010000: out_v[228] = 10'b0011001101;
    16'b0000010000001000: out_v[228] = 10'b1101000011;
    16'b0010000000011000: out_v[228] = 10'b1110111001;
    16'b0010001000000000: out_v[228] = 10'b1000100011;
    16'b0000011000011100: out_v[228] = 10'b0010111010;
    16'b0000000000010000: out_v[228] = 10'b0000011011;
    16'b0000001000000000: out_v[228] = 10'b1100100001;
    16'b0000000100001100: out_v[228] = 10'b0001011001;
    16'b0000010100000100: out_v[228] = 10'b0010001111;
    16'b0000010100001100: out_v[228] = 10'b1001010001;
    16'b0000010100011000: out_v[228] = 10'b0101111000;
    16'b0000001000111000: out_v[228] = 10'b1011011011;
    16'b0000010000001100: out_v[228] = 10'b1111000100;
    16'b0000000100000100: out_v[228] = 10'b0110001110;
    16'b0010001000011000: out_v[228] = 10'b0110110100;
    16'b0000010100000000: out_v[228] = 10'b0011000111;
    16'b0000010000000000: out_v[228] = 10'b1100110000;
    16'b0000000100000000: out_v[228] = 10'b0111100100;
    16'b0000000000000000: out_v[228] = 10'b0001101110;
    16'b0000010000100000: out_v[228] = 10'b1100100101;
    16'b0000000000100000: out_v[228] = 10'b1011001011;
    16'b0000010000000100: out_v[228] = 10'b0110100100;
    16'b0000010110100000: out_v[228] = 10'b1110100101;
    16'b0000010110100100: out_v[228] = 10'b0100101010;
    16'b0000010000100100: out_v[228] = 10'b1100010101;
    16'b0000010100100000: out_v[228] = 10'b1000101010;
    16'b0000010010100100: out_v[228] = 10'b0111011001;
    16'b0000010000010100: out_v[228] = 10'b1001011110;
    16'b0000010100100100: out_v[228] = 10'b1000100110;
    16'b0010010100100100: out_v[228] = 10'b1010011011;
    16'b0000000100100100: out_v[228] = 10'b1100000110;
    16'b0000000110100100: out_v[228] = 10'b1110100101;
    16'b0010010000000100: out_v[228] = 10'b1001111101;
    16'b0010010100000100: out_v[228] = 10'b0001100111;
    16'b0010010100100101: out_v[228] = 10'b0011001011;
    16'b0000010100100101: out_v[228] = 10'b1001111001;
    16'b0000000110100000: out_v[228] = 10'b1110110110;
    16'b0000000100100000: out_v[228] = 10'b1100100101;
    16'b0000010010100000: out_v[228] = 10'b0110100100;
    16'b0000011100010100: out_v[228] = 10'b0111001110;
    16'b0000010100010100: out_v[228] = 10'b1011001011;
    16'b0000000000000100: out_v[228] = 10'b1110101010;
    16'b0000000000101000: out_v[228] = 10'b0011001101;
    16'b0010000000000000: out_v[228] = 10'b1011100111;
    16'b0000000000101100: out_v[228] = 10'b0001110110;
    16'b0010000000001000: out_v[228] = 10'b0001001001;
    16'b0010000000000100: out_v[228] = 10'b0101100110;
    16'b0010000100000100: out_v[228] = 10'b0011001011;
    16'b0010000000011100: out_v[228] = 10'b0001010110;
    16'b0010000000001100: out_v[228] = 10'b0110011011;
    16'b0010000100000000: out_v[228] = 10'b0101011001;
    16'b0010000000101100: out_v[228] = 10'b1001111111;
    16'b0000000000111100: out_v[228] = 10'b0111100101;
    16'b0000000000100100: out_v[228] = 10'b1010100110;
    16'b0000010000101100: out_v[228] = 10'b1111101001;
    16'b0000000100001000: out_v[228] = 10'b1000011010;
    16'b0000000000010100: out_v[228] = 10'b0111101101;
    16'b0010001100011100: out_v[228] = 10'b1111000110;
    16'b0010001100010100: out_v[228] = 10'b1011001110;
    16'b0000010100001000: out_v[228] = 10'b1001110000;
    16'b0000001000010100: out_v[228] = 10'b0111111111;
    16'b0000011100011100: out_v[228] = 10'b0100010101;
    16'b0000001100010100: out_v[228] = 10'b1100100010;
    16'b0010000100011100: out_v[228] = 10'b1111000011;
    16'b0010001100010101: out_v[228] = 10'b1011101100;
    16'b0010001100011101: out_v[228] = 10'b0010011111;
    16'b0000001100000100: out_v[228] = 10'b1100110011;
    16'b0000000100010100: out_v[228] = 10'b0001011000;
    16'b0000001100011100: out_v[228] = 10'b1101000100;
    16'b0010001100000100: out_v[228] = 10'b1100110011;
    16'b0010001100000101: out_v[228] = 10'b1000010010;
    16'b0000001100011000: out_v[228] = 10'b0010100111;
    16'b0010001000011101: out_v[228] = 10'b0001110110;
    16'b0010001000011100: out_v[228] = 10'b0011110111;
    16'b0000001100010000: out_v[228] = 10'b1100011101;
    16'b0010000100011000: out_v[228] = 10'b1111110011;
    16'b0000011110111100: out_v[228] = 10'b0001001110;
    16'b0000010010011100: out_v[228] = 10'b0101001110;
    16'b0000010110111000: out_v[228] = 10'b1011001011;
    16'b0000010110111100: out_v[228] = 10'b1000001011;
    16'b0000011010110100: out_v[228] = 10'b1010001011;
    16'b0000010110101100: out_v[228] = 10'b0011001011;
    16'b0000010110011100: out_v[228] = 10'b1111100111;
    16'b0000011010111100: out_v[228] = 10'b1110100111;
    16'b0000011000010100: out_v[228] = 10'b1001000111;
    16'b0000010100111100: out_v[228] = 10'b1101001011;
    16'b0000010010111100: out_v[228] = 10'b1111101110;
    16'b0000011110110100: out_v[228] = 10'b0011101111;
    16'b0010001000010100: out_v[228] = 10'b0010001011;
    16'b0000001000000100: out_v[228] = 10'b1101111010;
    16'b0000011000000100: out_v[228] = 10'b0011100000;
    16'b1000001000010100: out_v[228] = 10'b1011011101;
    16'b0000010000010000: out_v[228] = 10'b1001110011;
    16'b0010010000011000: out_v[228] = 10'b1111100011;
    16'b0010011100011100: out_v[228] = 10'b0110100010;
    16'b0000000100010000: out_v[228] = 10'b0110001101;
    default: out_v[228] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100000100000001: out_v[229] = 10'b1100100001;
    16'b0000000100000001: out_v[229] = 10'b0001100100;
    16'b0110000100000001: out_v[229] = 10'b1000100100;
    16'b0110000100000000: out_v[229] = 10'b1010101011;
    16'b1100000100000001: out_v[229] = 10'b0101101001;
    16'b0101000100000000: out_v[229] = 10'b1001011011;
    16'b1110000100000001: out_v[229] = 10'b0000111011;
    16'b0010000100000000: out_v[229] = 10'b0000001011;
    16'b0100000000000000: out_v[229] = 10'b0001000111;
    16'b0101000000000000: out_v[229] = 10'b0001010011;
    16'b0010000100000001: out_v[229] = 10'b1101100001;
    16'b0100000100000000: out_v[229] = 10'b0100111001;
    16'b0110000000000000: out_v[229] = 10'b1100111010;
    16'b0101000100000001: out_v[229] = 10'b0000011101;
    16'b0100000000000001: out_v[229] = 10'b1100110110;
    16'b1010000100000001: out_v[229] = 10'b0111110010;
    16'b0010000000000000: out_v[229] = 10'b1010010100;
    16'b0111000100000001: out_v[229] = 10'b0011001001;
    16'b0000000100000000: out_v[229] = 10'b1110001000;
    16'b1110000000000001: out_v[229] = 10'b0011101110;
    16'b1110000100000000: out_v[229] = 10'b1011101100;
    16'b1000000100000001: out_v[229] = 10'b1001010010;
    16'b0111000100000000: out_v[229] = 10'b0000111111;
    16'b0000000000000000: out_v[229] = 10'b1001010110;
    16'b1000000000000000: out_v[229] = 10'b0011111100;
    16'b1000000100000000: out_v[229] = 10'b1111001010;
    16'b1100000000000000: out_v[229] = 10'b0001100110;
    16'b1100000100000000: out_v[229] = 10'b0111001110;
    16'b1110000000000000: out_v[229] = 10'b0000101110;
    16'b1101000000000000: out_v[229] = 10'b1001011110;
    16'b1111000100000000: out_v[229] = 10'b1101000111;
    16'b1100000000000001: out_v[229] = 10'b0110001111;
    16'b1101000100000001: out_v[229] = 10'b1101001111;
    16'b1101000100000000: out_v[229] = 10'b1101001000;
    16'b1111000000000000: out_v[229] = 10'b0010100101;
    16'b1010000000000000: out_v[229] = 10'b1101000100;
    16'b1010000100000000: out_v[229] = 10'b0100001100;
    16'b1001000100000000: out_v[229] = 10'b0110100111;
    16'b1000000000000001: out_v[229] = 10'b0100011100;
    16'b0000000000000001: out_v[229] = 10'b0110110001;
    16'b0010000000000001: out_v[229] = 10'b0111001110;
    16'b1010000000000001: out_v[229] = 10'b1010011011;
    16'b0110000000000001: out_v[229] = 10'b0000001001;
    16'b1001000000000000: out_v[229] = 10'b0111011010;
    16'b1001000100000001: out_v[229] = 10'b0010011010;
    16'b0001000000000000: out_v[229] = 10'b0011000011;
    16'b1000010100000000: out_v[229] = 10'b0111011000;
    16'b1000000100000101: out_v[229] = 10'b1000100011;
    16'b1000010100000001: out_v[229] = 10'b1100001110;
    16'b1000000100000010: out_v[229] = 10'b1011001101;
    16'b0000000100000010: out_v[229] = 10'b1111111010;
    16'b1000000100000100: out_v[229] = 10'b1010000010;
    16'b1100010100000000: out_v[229] = 10'b1101110001;
    default: out_v[229] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000010101000010: out_v[230] = 10'b0100101010;
    16'b0000000111000010: out_v[230] = 10'b1111001001;
    16'b0000000111100010: out_v[230] = 10'b1000001001;
    16'b0000000101100010: out_v[230] = 10'b0000111001;
    16'b0000000001000010: out_v[230] = 10'b1010001101;
    16'b0000010101000000: out_v[230] = 10'b1001000111;
    16'b0000000011100010: out_v[230] = 10'b0001111010;
    16'b0100010101000001: out_v[230] = 10'b1100001001;
    16'b0000000001100010: out_v[230] = 10'b1100101111;
    16'b0000010111000010: out_v[230] = 10'b1001011111;
    16'b0000000101000010: out_v[230] = 10'b1010110110;
    16'b0000000100100000: out_v[230] = 10'b0000101101;
    16'b1000000111100010: out_v[230] = 10'b0010101001;
    16'b0000000110000000: out_v[230] = 10'b0010110101;
    16'b0100010100000001: out_v[230] = 10'b1011101001;
    16'b0000010111100010: out_v[230] = 10'b1110001000;
    16'b0000010001000000: out_v[230] = 10'b0010011011;
    16'b0000000111100011: out_v[230] = 10'b0001000111;
    16'b0000010111100011: out_v[230] = 10'b1111001011;
    16'b0000000100100010: out_v[230] = 10'b1011001011;
    16'b0100010101000000: out_v[230] = 10'b1001010010;
    16'b0000010101100010: out_v[230] = 10'b1000100010;
    16'b0000000111000000: out_v[230] = 10'b0001011001;
    16'b0100000111100011: out_v[230] = 10'b1111100000;
    16'b0000000101000000: out_v[230] = 10'b0011011001;
    16'b0000000001000000: out_v[230] = 10'b0000111001;
    16'b1000000101100010: out_v[230] = 10'b1011101010;
    16'b0000010111000000: out_v[230] = 10'b1000001111;
    16'b0100000110000001: out_v[230] = 10'b1010110010;
    16'b0000000100000000: out_v[230] = 10'b1010100001;
    16'b0000010001000010: out_v[230] = 10'b1011101010;
    16'b0000000101100011: out_v[230] = 10'b0110110111;
    16'b0100010111000001: out_v[230] = 10'b0000011110;
    16'b0100010110000001: out_v[230] = 10'b1011000111;
    16'b0000010111000011: out_v[230] = 10'b0110001001;
    16'b0100010111100011: out_v[230] = 10'b0100001001;
    16'b0100010111000000: out_v[230] = 10'b0111110001;
    16'b0000000110000001: out_v[230] = 10'b0010100010;
    16'b0100000001000000: out_v[230] = 10'b0100100110;
    16'b0100000001000001: out_v[230] = 10'b0001001110;
    16'b0100000000000001: out_v[230] = 10'b1101010100;
    16'b0000000100000001: out_v[230] = 10'b1111011001;
    16'b0100000000000010: out_v[230] = 10'b0001000011;
    16'b0100000000000000: out_v[230] = 10'b0110100111;
    16'b0100000111000001: out_v[230] = 10'b0011111010;
    16'b0000000000000001: out_v[230] = 10'b1000110100;
    16'b0000000101000001: out_v[230] = 10'b0100001000;
    16'b0100000101000001: out_v[230] = 10'b0011011101;
    16'b0000000010000001: out_v[230] = 10'b0001111011;
    16'b0000000111000001: out_v[230] = 10'b1110010011;
    16'b0100000001000011: out_v[230] = 10'b1010100010;
    16'b0000000000000010: out_v[230] = 10'b1101011010;
    16'b0100000000000011: out_v[230] = 10'b1010111111;
    16'b0000000001000001: out_v[230] = 10'b0101100100;
    16'b0100000101000000: out_v[230] = 10'b1001000010;
    16'b0100000100000001: out_v[230] = 10'b1110100001;
    16'b0100000001000010: out_v[230] = 10'b0011000110;
    16'b0000000111000011: out_v[230] = 10'b1100110100;
    16'b0100010010000001: out_v[230] = 10'b1100101011;
    16'b0100000110100011: out_v[230] = 10'b1010010100;
    16'b0100010110100001: out_v[230] = 10'b0000111010;
    16'b0100010000100001: out_v[230] = 10'b1001010010;
    16'b0100010110100011: out_v[230] = 10'b1100010100;
    16'b0100010100100001: out_v[230] = 10'b0011001011;
    16'b0100010000000011: out_v[230] = 10'b0000111000;
    16'b1100010000000011: out_v[230] = 10'b1111100111;
    16'b0100010100100011: out_v[230] = 10'b1001110110;
    16'b0100000110100001: out_v[230] = 10'b1110000100;
    16'b0101010110100001: out_v[230] = 10'b0111101110;
    16'b0100010100000011: out_v[230] = 10'b1101000100;
    16'b1100010111000011: out_v[230] = 10'b0011110100;
    16'b0100000000100001: out_v[230] = 10'b1000010110;
    16'b0100010111100001: out_v[230] = 10'b0001110110;
    16'b1100010110000011: out_v[230] = 10'b0100110110;
    16'b0100000110000011: out_v[230] = 10'b1010111101;
    16'b0100010000100011: out_v[230] = 10'b0001000000;
    16'b0100000100100001: out_v[230] = 10'b1110011111;
    16'b1100000110000011: out_v[230] = 10'b0111000110;
    16'b0000000000100001: out_v[230] = 10'b1110000110;
    16'b0100010000000001: out_v[230] = 10'b0001000111;
    16'b1100010111100011: out_v[230] = 10'b0000100111;
    16'b1000000111000011: out_v[230] = 10'b1011111111;
    16'b0000000110100011: out_v[230] = 10'b0010101101;
    16'b0100010101100001: out_v[230] = 10'b0111000110;
    16'b0000000110100001: out_v[230] = 10'b1001000101;
    16'b0100010110000011: out_v[230] = 10'b1001101110;
    16'b0000010000000001: out_v[230] = 10'b0000001111;
    16'b0100010111000011: out_v[230] = 10'b0100111011;
    16'b1100010100000011: out_v[230] = 10'b1001101001;
    16'b0100010010100001: out_v[230] = 10'b1101100110;
    16'b0000010100100001: out_v[230] = 10'b1011000110;
    16'b0000010011000000: out_v[230] = 10'b1100101011;
    16'b0000010001100010: out_v[230] = 10'b0100101100;
    16'b0000000011000010: out_v[230] = 10'b1011101101;
    16'b0000010000000010: out_v[230] = 10'b0110010001;
    16'b0000010011000010: out_v[230] = 10'b0100101110;
    16'b1000010001100010: out_v[230] = 10'b0010101101;
    16'b1000010111100010: out_v[230] = 10'b0010011111;
    16'b0000010011100010: out_v[230] = 10'b1100011111;
    16'b0000010100000000: out_v[230] = 10'b1101000010;
    16'b0000010110100010: out_v[230] = 10'b0011011111;
    16'b0000010000100010: out_v[230] = 10'b0111110000;
    16'b0000000110000010: out_v[230] = 10'b0000011110;
    16'b0000010110000011: out_v[230] = 10'b1001110011;
    16'b0000010000000011: out_v[230] = 10'b0110000010;
    16'b0100010001001000: out_v[230] = 10'b0011110101;
    16'b0000010110000010: out_v[230] = 10'b0010010010;
    16'b0100010011000001: out_v[230] = 10'b0111111000;
    16'b0100010001000000: out_v[230] = 10'b0011110001;
    16'b0100010000000000: out_v[230] = 10'b0110010100;
    16'b0100010001000001: out_v[230] = 10'b0100110000;
    16'b0000010010000000: out_v[230] = 10'b0010000011;
    16'b0100010001001001: out_v[230] = 10'b0000111100;
    16'b0000010000000000: out_v[230] = 10'b0101011000;
    16'b0100000111000000: out_v[230] = 10'b1010011101;
    16'b1000010000100000: out_v[230] = 10'b1001110111;
    16'b0100010011000000: out_v[230] = 10'b0111010011;
    16'b0000010010000010: out_v[230] = 10'b1010100010;
    16'b1000010110100000: out_v[230] = 10'b0111011011;
    16'b0000010110000001: out_v[230] = 10'b0110010000;
    16'b0000010110000000: out_v[230] = 10'b0101010011;
    16'b0100010110000010: out_v[230] = 10'b0011010011;
    16'b0000010001001000: out_v[230] = 10'b0101010011;
    16'b1000010110100010: out_v[230] = 10'b1011011101;
    16'b0000010100000010: out_v[230] = 10'b1100001100;
    16'b0100000010000000: out_v[230] = 10'b0111111000;
    16'b0100000010000001: out_v[230] = 10'b0011101000;
    16'b0100000101000010: out_v[230] = 10'b1011110111;
    16'b0000010100100010: out_v[230] = 10'b1111001001;
    16'b0000000000000000: out_v[230] = 10'b1110001101;
    16'b0000000010000000: out_v[230] = 10'b1100100101;
    16'b0100000101000011: out_v[230] = 10'b1000111011;
    16'b0100000011000000: out_v[230] = 10'b1000001100;
    16'b0000000100000010: out_v[230] = 10'b0001101101;
    16'b1000010101100010: out_v[230] = 10'b1011100101;
    16'b0000000011000000: out_v[230] = 10'b0111101000;
    16'b0000000100001010: out_v[230] = 10'b0111100110;
    16'b0100000011000001: out_v[230] = 10'b1111100000;
    16'b0000010001100011: out_v[230] = 10'b0011011000;
    16'b0100010101100011: out_v[230] = 10'b1001100000;
    16'b0100000000100011: out_v[230] = 10'b0101000000;
    16'b0000000000100011: out_v[230] = 10'b0111000101;
    16'b0000010000100011: out_v[230] = 10'b0000111011;
    16'b0000000001000011: out_v[230] = 10'b1111001100;
    16'b0100010001100011: out_v[230] = 10'b0011101011;
    16'b0000010000100001: out_v[230] = 10'b0111111001;
    16'b0000010101000001: out_v[230] = 10'b1001100111;
    16'b0000010101100011: out_v[230] = 10'b0101100000;
    16'b0000010001000011: out_v[230] = 10'b1001100110;
    16'b0000010100000001: out_v[230] = 10'b1100100000;
    16'b0100010001000011: out_v[230] = 10'b0101100011;
    16'b0000010001000001: out_v[230] = 10'b1101001000;
    16'b0000000000000011: out_v[230] = 10'b1111100111;
    16'b0000000001100011: out_v[230] = 10'b1011000101;
    16'b0000010101000011: out_v[230] = 10'b1110010001;
    16'b0100010000100010: out_v[230] = 10'b1111101111;
    16'b0100010111001001: out_v[230] = 10'b0011101010;
    16'b0100010111001000: out_v[230] = 10'b0111100111;
    16'b0100010011001001: out_v[230] = 10'b0111101111;
    16'b0000010111001010: out_v[230] = 10'b0001111111;
    16'b0000010011001010: out_v[230] = 10'b1111000110;
    16'b0100010011001000: out_v[230] = 10'b1000000110;
    16'b0100010010000000: out_v[230] = 10'b0010000101;
    16'b0000010011001000: out_v[230] = 10'b0111100001;
    16'b0000010111001000: out_v[230] = 10'b1101010010;
    16'b0100010111001010: out_v[230] = 10'b1011010011;
    16'b0000010010000110: out_v[230] = 10'b1011010111;
    16'b0100010101001000: out_v[230] = 10'b1001001111;
    16'b0100000111001001: out_v[230] = 10'b0011000011;
    16'b0100000111001000: out_v[230] = 10'b0110110001;
    16'b0100010101001001: out_v[230] = 10'b1100000010;
    16'b0100000011001000: out_v[230] = 10'b0111101010;
    16'b0000010101001000: out_v[230] = 10'b1000000100;
    16'b0000010010000001: out_v[230] = 10'b0111011010;
    16'b0000000101000011: out_v[230] = 10'b1111110101;
    16'b0100000111000011: out_v[230] = 10'b0101100110;
    16'b0100010101000011: out_v[230] = 10'b1101011011;
    16'b0000000100000011: out_v[230] = 10'b1101011011;
    16'b0000000110000011: out_v[230] = 10'b0100001101;
    16'b0000000011000011: out_v[230] = 10'b1100011001;
    16'b0100010100000000: out_v[230] = 10'b1101001001;
    16'b0000010100000011: out_v[230] = 10'b1110000101;
    16'b0000010010000011: out_v[230] = 10'b1101110010;
    16'b1000010010100000: out_v[230] = 10'b1001010110;
    16'b0100000101001000: out_v[230] = 10'b1001001101;
    16'b0000000010000010: out_v[230] = 10'b1010101110;
    default: out_v[230] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1011000000000000: out_v[231] = 10'b1010001001;
    16'b0011000000000000: out_v[231] = 10'b1000101001;
    16'b0001000000000010: out_v[231] = 10'b0010011101;
    16'b0010000000000000: out_v[231] = 10'b1100011001;
    16'b0000000000000000: out_v[231] = 10'b1010101001;
    16'b0001000000000000: out_v[231] = 10'b1001100101;
    16'b1010000000000000: out_v[231] = 10'b0101101011;
    16'b0011000100000000: out_v[231] = 10'b0010010100;
    16'b0011000000000010: out_v[231] = 10'b1001100110;
    16'b1011000100000000: out_v[231] = 10'b0011011101;
    16'b1000000000000000: out_v[231] = 10'b0100110111;
    16'b1001000000000000: out_v[231] = 10'b1111011000;
    16'b0011000000010000: out_v[231] = 10'b1001011100;
    16'b0001000100000010: out_v[231] = 10'b0100101011;
    16'b1000000000000010: out_v[231] = 10'b0000111011;
    16'b1001000000000010: out_v[231] = 10'b1111110000;
    16'b0010000000010000: out_v[231] = 10'b0010010100;
    16'b0000000000010000: out_v[231] = 10'b1110111001;
    16'b0001000100000000: out_v[231] = 10'b1101110001;
    16'b1000000000010000: out_v[231] = 10'b0001011110;
    16'b1001000000010000: out_v[231] = 10'b1100101010;
    16'b0001000000010000: out_v[231] = 10'b1000000110;
    16'b0001000000010010: out_v[231] = 10'b0001010101;
    16'b0001000100010000: out_v[231] = 10'b0101010110;
    16'b0000000000010010: out_v[231] = 10'b1010011101;
    16'b0010000000010010: out_v[231] = 10'b1011101110;
    16'b0011000000010010: out_v[231] = 10'b1011011010;
    16'b1011000000010000: out_v[231] = 10'b0110111010;
    16'b1010000000010000: out_v[231] = 10'b0110011100;
    16'b0011000000001000: out_v[231] = 10'b1101101101;
    16'b0000100000010100: out_v[231] = 10'b0101001111;
    16'b0011000100010000: out_v[231] = 10'b1000011110;
    16'b0010000100010000: out_v[231] = 10'b1000010000;
    16'b1011000100010000: out_v[231] = 10'b1001010001;
    16'b0000000000010100: out_v[231] = 10'b0001111101;
    16'b0001000000010100: out_v[231] = 10'b1000111010;
    16'b0000000000000100: out_v[231] = 10'b0001111010;
    16'b0001100000010100: out_v[231] = 10'b0010010001;
    16'b0000100000000100: out_v[231] = 10'b1010010100;
    16'b1001100000010100: out_v[231] = 10'b1011101010;
    16'b0001100000000100: out_v[231] = 10'b1000110010;
    16'b0001000000000100: out_v[231] = 10'b0010110101;
    16'b0011000001010000: out_v[231] = 10'b1101011001;
    16'b0011000001000000: out_v[231] = 10'b1111100110;
    16'b0001000001010000: out_v[231] = 10'b1010000111;
    16'b0010000001010000: out_v[231] = 10'b1111100111;
    16'b0010000100000000: out_v[231] = 10'b1110010000;
    16'b0000000100010000: out_v[231] = 10'b0101110011;
    16'b1001000100010000: out_v[231] = 10'b0101111110;
    16'b1001000100000000: out_v[231] = 10'b1000001001;
    16'b0000000100000000: out_v[231] = 10'b1011100010;
    default: out_v[231] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000000011100: out_v[232] = 10'b0010011011;
    16'b0000011000011101: out_v[232] = 10'b1111010111;
    16'b0000010000011101: out_v[232] = 10'b0010110000;
    16'b0000000000001101: out_v[232] = 10'b0011101000;
    16'b0000110000011101: out_v[232] = 10'b0000110011;
    16'b0000010000001001: out_v[232] = 10'b0101011101;
    16'b0000010000001000: out_v[232] = 10'b1001001010;
    16'b0000010000001101: out_v[232] = 10'b1001001000;
    16'b0000010000000101: out_v[232] = 10'b1001001111;
    16'b0000100000011101: out_v[232] = 10'b0010110011;
    16'b0010010000001101: out_v[232] = 10'b0101011100;
    16'b0010110000111101: out_v[232] = 10'b0001011010;
    16'b0000010000001100: out_v[232] = 10'b1111100100;
    16'b0000000000011101: out_v[232] = 10'b0010110101;
    16'b0000010000010101: out_v[232] = 10'b0010110001;
    16'b0000010000000100: out_v[232] = 10'b1100011110;
    16'b0000000000010101: out_v[232] = 10'b0010001111;
    16'b0000011000001101: out_v[232] = 10'b0111011011;
    16'b0010010000101101: out_v[232] = 10'b0110110101;
    16'b0000000000000101: out_v[232] = 10'b0111001111;
    16'b0010100000111101: out_v[232] = 10'b1110001010;
    16'b0000010000011001: out_v[232] = 10'b1111110011;
    16'b0000110000001101: out_v[232] = 10'b1010111001;
    16'b0010000000011101: out_v[232] = 10'b0011101001;
    16'b0000010000011100: out_v[232] = 10'b0011111110;
    16'b0000010000000000: out_v[232] = 10'b0001011101;
    16'b0000010000000001: out_v[232] = 10'b1001101101;
    16'b0000000000000100: out_v[232] = 10'b1001111101;
    16'b0000000000001100: out_v[232] = 10'b1000101110;
    16'b0010010000111101: out_v[232] = 10'b1111000110;
    16'b0010110000110000: out_v[232] = 10'b0010100101;
    16'b0010000000111101: out_v[232] = 10'b1000110011;
    16'b0010000000010101: out_v[232] = 10'b1100101011;
    16'b0000110000011001: out_v[232] = 10'b1010101101;
    16'b0010110000111001: out_v[232] = 10'b0111011011;
    16'b0000110000111101: out_v[232] = 10'b0010001000;
    16'b0010100000110000: out_v[232] = 10'b1011100011;
    16'b0010100000100101: out_v[232] = 10'b1010101010;
    16'b0010000000100001: out_v[232] = 10'b1001010000;
    16'b0010000000100101: out_v[232] = 10'b0011110011;
    16'b0010100000100000: out_v[232] = 10'b0111011100;
    16'b0000100000100101: out_v[232] = 10'b0000110010;
    16'b0010101000110000: out_v[232] = 10'b1001001110;
    16'b0010100000110001: out_v[232] = 10'b1101001000;
    16'b0010100000100001: out_v[232] = 10'b0111111100;
    16'b0010000000100000: out_v[232] = 10'b1011100110;
    16'b0000100000010000: out_v[232] = 10'b0000111110;
    16'b0000100000100001: out_v[232] = 10'b1100011001;
    16'b0000100000100000: out_v[232] = 10'b1110010010;
    16'b0010000000100100: out_v[232] = 10'b0100001011;
    16'b0000000000100101: out_v[232] = 10'b1100011011;
    16'b0010100000110101: out_v[232] = 10'b1000001010;
    16'b0000100000110000: out_v[232] = 10'b1110101000;
    16'b0000100000010101: out_v[232] = 10'b0111100110;
    16'b0000000000000000: out_v[232] = 10'b1100100111;
    16'b0000100000011000: out_v[232] = 10'b0011111000;
    16'b0000010000011000: out_v[232] = 10'b1100001010;
    16'b0010100000110111: out_v[232] = 10'b0111011110;
    16'b0000010000010000: out_v[232] = 10'b0010000111;
    16'b0010100000111000: out_v[232] = 10'b1000001011;
    16'b0000000000010001: out_v[232] = 10'b0000101111;
    16'b0000000000011001: out_v[232] = 10'b0010010100;
    16'b0000110000011000: out_v[232] = 10'b1000011010;
    16'b0000000000010000: out_v[232] = 10'b1010101101;
    16'b0000100000011001: out_v[232] = 10'b0110110000;
    16'b0000110000010000: out_v[232] = 10'b1110100010;
    16'b0000010000011010: out_v[232] = 10'b1110101110;
    16'b0000100000010001: out_v[232] = 10'b0111101111;
    16'b0010100000101000: out_v[232] = 10'b1000011111;
    16'b0010110000111000: out_v[232] = 10'b1101000110;
    16'b0010100000111001: out_v[232] = 10'b1011001100;
    16'b0000100000010111: out_v[232] = 10'b0100011101;
    16'b0010010000011000: out_v[232] = 10'b1000110011;
    16'b0000010000010001: out_v[232] = 10'b1011001010;
    16'b0010110000101000: out_v[232] = 10'b1011011100;
    16'b0010010000001000: out_v[232] = 10'b0101101110;
    16'b0000000000011000: out_v[232] = 10'b0010011100;
    16'b0010000000101000: out_v[232] = 10'b0010101111;
    16'b0010100000010101: out_v[232] = 10'b1111100001;
    16'b0010110000011000: out_v[232] = 10'b1011000101;
    16'b0010100000101100: out_v[232] = 10'b0110101011;
    16'b0010100000101101: out_v[232] = 10'b0011110000;
    16'b0010100100111101: out_v[232] = 10'b0001110100;
    16'b0010100100101101: out_v[232] = 10'b1001001000;
    16'b0010101000111100: out_v[232] = 10'b0111001011;
    16'b0010000000101101: out_v[232] = 10'b0110111001;
    16'b0010101000111101: out_v[232] = 10'b0011001011;
    16'b0010100000110100: out_v[232] = 10'b0110011110;
    16'b0010100000111100: out_v[232] = 10'b1101000010;
    16'b0010100100111100: out_v[232] = 10'b1010111111;
    16'b0010110000110101: out_v[232] = 10'b1111000010;
    16'b0010101000110101: out_v[232] = 10'b0000011110;
    16'b0010101000110001: out_v[232] = 10'b1111000101;
    16'b0010000000101100: out_v[232] = 10'b0111001101;
    16'b0010100000100100: out_v[232] = 10'b1100011101;
    16'b0000100000101101: out_v[232] = 10'b0101011010;
    16'b0010100100110101: out_v[232] = 10'b1001101001;
    16'b0010101000101101: out_v[232] = 10'b0111110111;
    16'b0010101010111101: out_v[232] = 10'b0000011011;
    16'b0010000000010001: out_v[232] = 10'b1000101111;
    16'b0000100000000000: out_v[232] = 10'b1110011010;
    16'b0010100000010001: out_v[232] = 10'b0111100111;
    16'b0010100000010000: out_v[232] = 10'b0110100001;
    16'b0010100000010100: out_v[232] = 10'b1100000000;
    16'b0010110000010101: out_v[232] = 10'b1001110111;
    16'b0000000000001000: out_v[232] = 10'b1001110000;
    16'b0000100000010100: out_v[232] = 10'b1111110110;
    16'b0000110000010001: out_v[232] = 10'b1111100010;
    16'b0010100000011000: out_v[232] = 10'b0110010111;
    16'b0010000000010000: out_v[232] = 10'b1001010010;
    16'b0000000000010100: out_v[232] = 10'b0001011111;
    16'b0000000000000001: out_v[232] = 10'b1101011010;
    16'b0000100000000100: out_v[232] = 10'b1100010101;
    16'b0010000000011000: out_v[232] = 10'b1000011001;
    16'b0000110000010101: out_v[232] = 10'b0000110110;
    16'b0010000000110101: out_v[232] = 10'b0101110010;
    16'b0000010000010100: out_v[232] = 10'b0101011001;
    16'b0000100000000101: out_v[232] = 10'b0100101100;
    16'b0010010000010101: out_v[232] = 10'b1001011011;
    16'b0010000000000101: out_v[232] = 10'b1001101011;
    16'b0010001000101101: out_v[232] = 10'b1111011101;
    16'b0010001000000101: out_v[232] = 10'b0011011111;
    16'b0010000000001101: out_v[232] = 10'b1010111010;
    16'b0010000000001100: out_v[232] = 10'b0001101110;
    16'b0000001000000101: out_v[232] = 10'b1000010101;
    16'b0010000000000000: out_v[232] = 10'b1101100110;
    16'b0010001000100101: out_v[232] = 10'b1011100011;
    16'b0010000000000001: out_v[232] = 10'b1110001000;
    16'b0010010000100101: out_v[232] = 10'b0100110000;
    16'b0010110000101101: out_v[232] = 10'b0001100001;
    16'b0010001000001101: out_v[232] = 10'b1110011111;
    16'b0010000000000100: out_v[232] = 10'b0111111011;
    16'b0000000000001001: out_v[232] = 10'b0110101100;
    16'b0010000000001001: out_v[232] = 10'b0110011001;
    16'b1000000000001001: out_v[232] = 10'b1110110010;
    16'b0010000000101001: out_v[232] = 10'b1101100111;
    16'b1010100000111001: out_v[232] = 10'b1111111010;
    16'b1000000000001000: out_v[232] = 10'b1111001111;
    16'b0010000000001000: out_v[232] = 10'b1100101001;
    16'b0010010000001001: out_v[232] = 10'b1101001010;
    16'b0010100000101001: out_v[232] = 10'b1110100001;
    16'b1000000000000001: out_v[232] = 10'b0011001100;
    16'b1000100000011001: out_v[232] = 10'b1101000011;
    16'b0010010000101001: out_v[232] = 10'b0010100111;
    16'b0000101000010001: out_v[232] = 10'b0111110011;
    16'b0000100000110101: out_v[232] = 10'b0111100100;
    16'b0000001000010001: out_v[232] = 10'b1110000111;
    16'b0000100000111101: out_v[232] = 10'b1011000001;
    16'b0000001000010000: out_v[232] = 10'b0110011000;
    16'b0000100000110001: out_v[232] = 10'b1110101000;
    16'b0000101000010000: out_v[232] = 10'b0011010000;
    16'b0000100000011100: out_v[232] = 10'b0100010011;
    16'b0000001000000000: out_v[232] = 10'b0111001100;
    16'b0010000000010100: out_v[232] = 10'b0100110111;
    16'b0010100000011101: out_v[232] = 10'b0100101001;
    16'b0010001000010101: out_v[232] = 10'b0010111111;
    16'b0010101000010101: out_v[232] = 10'b0100011111;
    default: out_v[232] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1100000001000001: out_v[233] = 10'b0010100111;
    16'b1000110101000001: out_v[233] = 10'b0001101011;
    16'b1100110100100001: out_v[233] = 10'b1110000111;
    16'b1100110101100001: out_v[233] = 10'b0100010011;
    16'b1100110001100001: out_v[233] = 10'b1110100100;
    16'b1000110100000001: out_v[233] = 10'b1101010011;
    16'b0000110000100000: out_v[233] = 10'b1101011111;
    16'b0100110101100000: out_v[233] = 10'b0111010001;
    16'b1100111001100000: out_v[233] = 10'b1101101110;
    16'b1100000001000000: out_v[233] = 10'b0111010111;
    16'b1100110101000001: out_v[233] = 10'b1111111100;
    16'b1100100001000001: out_v[233] = 10'b0100011011;
    16'b0100110101100001: out_v[233] = 10'b0111011110;
    16'b1100100001100001: out_v[233] = 10'b1011011011;
    16'b1100111001100001: out_v[233] = 10'b0010111011;
    16'b0100110101000001: out_v[233] = 10'b0100000100;
    16'b1100111101100001: out_v[233] = 10'b1111011111;
    16'b0100100101000001: out_v[233] = 10'b0100000111;
    16'b1000000001000001: out_v[233] = 10'b1111000010;
    16'b1100110101100000: out_v[233] = 10'b0110011110;
    16'b1100110001100000: out_v[233] = 10'b0000100111;
    16'b1000110100100001: out_v[233] = 10'b1110111110;
    16'b1100111101100000: out_v[233] = 10'b0110011111;
    16'b1100010101100000: out_v[233] = 10'b0011111011;
    16'b1100001001000001: out_v[233] = 10'b0110001011;
    16'b1000110100100000: out_v[233] = 10'b0111111111;
    16'b0100010101100000: out_v[233] = 10'b1000000011;
    16'b1100100101000001: out_v[233] = 10'b1011000100;
    16'b1100110001000001: out_v[233] = 10'b0110011001;
    16'b1000110101100001: out_v[233] = 10'b1011001101;
    16'b1000100100000001: out_v[233] = 10'b1000000101;
    16'b1100101001100001: out_v[233] = 10'b0111001011;
    16'b1000100101000001: out_v[233] = 10'b1111111010;
    16'b0100000001000001: out_v[233] = 10'b1000101100;
    16'b1100010101100001: out_v[233] = 10'b1011011110;
    16'b1100101001000001: out_v[233] = 10'b0101110101;
    16'b1000110001100001: out_v[233] = 10'b0011111110;
    16'b1000110101100000: out_v[233] = 10'b1110111010;
    16'b0100111101100000: out_v[233] = 10'b1001111000;
    16'b1000000100000000: out_v[233] = 10'b0000101010;
    16'b1000000000000000: out_v[233] = 10'b1001001011;
    16'b0000000001000000: out_v[233] = 10'b1110110001;
    16'b0100000001000000: out_v[233] = 10'b1100000110;
    16'b1000000001000000: out_v[233] = 10'b0100110111;
    16'b0000000100000000: out_v[233] = 10'b0011100011;
    16'b0100000000000000: out_v[233] = 10'b0010111000;
    16'b0100001001000000: out_v[233] = 10'b0111110000;
    16'b0000000000000000: out_v[233] = 10'b1100110011;
    16'b0100001000000000: out_v[233] = 10'b1100001000;
    16'b1100001001000000: out_v[233] = 10'b0001010100;
    16'b1100001101000000: out_v[233] = 10'b0011100011;
    16'b1000001001000000: out_v[233] = 10'b0010011100;
    16'b1000100101000010: out_v[233] = 10'b1010011001;
    16'b1000001100000010: out_v[233] = 10'b1111010111;
    16'b0000100000000000: out_v[233] = 10'b1100101011;
    16'b0000101001000000: out_v[233] = 10'b1110101010;
    16'b1000100101000000: out_v[233] = 10'b1100011010;
    16'b1000000101000000: out_v[233] = 10'b0110111100;
    16'b0000100001000000: out_v[233] = 10'b0010011100;
    16'b1000000101000001: out_v[233] = 10'b1010011110;
    16'b0000001001000000: out_v[233] = 10'b0101101001;
    16'b0000100001100000: out_v[233] = 10'b1010111101;
    16'b1000101101000011: out_v[233] = 10'b1111111011;
    16'b1000001101000000: out_v[233] = 10'b0100110101;
    16'b1000101101000000: out_v[233] = 10'b1110000011;
    16'b1000001101000001: out_v[233] = 10'b0011110010;
    16'b0000100001000001: out_v[233] = 10'b1001100100;
    16'b1000101001000000: out_v[233] = 10'b1110001110;
    16'b1000101101000001: out_v[233] = 10'b0111110100;
    16'b0000100000100000: out_v[233] = 10'b0100000110;
    16'b1000100101000011: out_v[233] = 10'b1110100110;
    16'b0000000000100000: out_v[233] = 10'b1000000110;
    16'b0000100101000000: out_v[233] = 10'b0110010110;
    16'b0000000101000000: out_v[233] = 10'b0111110000;
    16'b0000101001100000: out_v[233] = 10'b1111101111;
    16'b1100001101000001: out_v[233] = 10'b1001100101;
    16'b1000001101100000: out_v[233] = 10'b1101110111;
    16'b1100000101000000: out_v[233] = 10'b1011001111;
    16'b1000001001100000: out_v[233] = 10'b1000010101;
    16'b0000110001000001: out_v[233] = 10'b0101100011;
    16'b0000110101000001: out_v[233] = 10'b0110000110;
    16'b0000100101000010: out_v[233] = 10'b0101111011;
    16'b0100000101000000: out_v[233] = 10'b0110111000;
    16'b0100001101000000: out_v[233] = 10'b0010111001;
    16'b1100000101000001: out_v[233] = 10'b0111110000;
    16'b1100001001100001: out_v[233] = 10'b1000111011;
    16'b0100001101100001: out_v[233] = 10'b1011100110;
    16'b0100001101000001: out_v[233] = 10'b0101001011;
    16'b1100001101100001: out_v[233] = 10'b0011001000;
    16'b0100001100000000: out_v[233] = 10'b1001001011;
    16'b1100001001100000: out_v[233] = 10'b1010101110;
    16'b0100001001100000: out_v[233] = 10'b1010101001;
    16'b0100000101100001: out_v[233] = 10'b0111111011;
    16'b0100000101000001: out_v[233] = 10'b1111011000;
    16'b0100000000000001: out_v[233] = 10'b0011110010;
    16'b1000100000000000: out_v[233] = 10'b0001111100;
    16'b0100100001100000: out_v[233] = 10'b0000111010;
    16'b0000000001000001: out_v[233] = 10'b0111110000;
    16'b1000010000000001: out_v[233] = 10'b0110011000;
    16'b0000100000100001: out_v[233] = 10'b1000101110;
    16'b1000000000000001: out_v[233] = 10'b0010000001;
    16'b0000000000000001: out_v[233] = 10'b0000111111;
    16'b0100001000000001: out_v[233] = 10'b0011011101;
    16'b0100010000000001: out_v[233] = 10'b0111011100;
    16'b1000100000000001: out_v[233] = 10'b1101110111;
    16'b0100100000100000: out_v[233] = 10'b0011111010;
    16'b0000010000000001: out_v[233] = 10'b0100001111;
    16'b0100100000000001: out_v[233] = 10'b1110010000;
    16'b0100000000100000: out_v[233] = 10'b0010011001;
    16'b0000110000000001: out_v[233] = 10'b1001011101;
    16'b0100110000000001: out_v[233] = 10'b0010001110;
    16'b0100100000000000: out_v[233] = 10'b1110111010;
    16'b0100100001000001: out_v[233] = 10'b1110100001;
    16'b0100100000100001: out_v[233] = 10'b1100111010;
    16'b0100100001000000: out_v[233] = 10'b1000110011;
    16'b0000100000000001: out_v[233] = 10'b1010010010;
    16'b0100101000000001: out_v[233] = 10'b0010011111;
    16'b0000110000100001: out_v[233] = 10'b0010110001;
    16'b1000100000100000: out_v[233] = 10'b1001110010;
    16'b1000010100000000: out_v[233] = 10'b0001110001;
    16'b1100100001000000: out_v[233] = 10'b1001111110;
    16'b0000110000000000: out_v[233] = 10'b0111100010;
    16'b0100000100000000: out_v[233] = 10'b1001001100;
    16'b1100000100000000: out_v[233] = 10'b1111000010;
    16'b1100000000000000: out_v[233] = 10'b0101001100;
    16'b1000100100000000: out_v[233] = 10'b1101000011;
    16'b0000010000000000: out_v[233] = 10'b1000101010;
    16'b1100000101100001: out_v[233] = 10'b0110100000;
    16'b1100000001100001: out_v[233] = 10'b1000111110;
    16'b0100000001000010: out_v[233] = 10'b1011000001;
    16'b1100100001100011: out_v[233] = 10'b1101011110;
    16'b1000000001000011: out_v[233] = 10'b1101110111;
    16'b0000001000100001: out_v[233] = 10'b0111100001;
    16'b1100000001000011: out_v[233] = 10'b0011010011;
    16'b1100000001000010: out_v[233] = 10'b1111010010;
    16'b1000100001100011: out_v[233] = 10'b0110110001;
    16'b0000000000100001: out_v[233] = 10'b1101000011;
    16'b1000000001000010: out_v[233] = 10'b0110111011;
    16'b0000100001100011: out_v[233] = 10'b1001101001;
    16'b1001000000000000: out_v[233] = 10'b0001001100;
    16'b1000110001100011: out_v[233] = 10'b1000110011;
    16'b0000011000100001: out_v[233] = 10'b0110101111;
    16'b0000111000100001: out_v[233] = 10'b1111100100;
    16'b0000000001000010: out_v[233] = 10'b1111010010;
    16'b1100000001100011: out_v[233] = 10'b0001011110;
    16'b0000001000000001: out_v[233] = 10'b0110100111;
    16'b1000100001000011: out_v[233] = 10'b1110001111;
    16'b1000111000100001: out_v[233] = 10'b1111101011;
    16'b0000000001100011: out_v[233] = 10'b1110001011;
    16'b1000000001100011: out_v[233] = 10'b0110110001;
    16'b1000100001100001: out_v[233] = 10'b1010110110;
    16'b0000000001000011: out_v[233] = 10'b1101101011;
    16'b1001100000000000: out_v[233] = 10'b1101010011;
    16'b1001100000000001: out_v[233] = 10'b0111111010;
    16'b0000101000100001: out_v[233] = 10'b1101101110;
    16'b0100000000000101: out_v[233] = 10'b0111110100;
    16'b1000010100000001: out_v[233] = 10'b0100000110;
    16'b0000000000000101: out_v[233] = 10'b1011100111;
    16'b0100000000000100: out_v[233] = 10'b0010011010;
    16'b0100010000000101: out_v[233] = 10'b0101010111;
    16'b1100011001000001: out_v[233] = 10'b0110000011;
    16'b1000010101000001: out_v[233] = 10'b1011111010;
    16'b0100010101000000: out_v[233] = 10'b0111011100;
    16'b0100100101000000: out_v[233] = 10'b0100111101;
    16'b0000010100000001: out_v[233] = 10'b1110010010;
    16'b0100010001000001: out_v[233] = 10'b1110000000;
    16'b0100010101000001: out_v[233] = 10'b1111011011;
    16'b1100001000000000: out_v[233] = 10'b1111100111;
    16'b1100010001000001: out_v[233] = 10'b0110110010;
    16'b1100010101000001: out_v[233] = 10'b1001011111;
    16'b1100010001000000: out_v[233] = 10'b1001110000;
    16'b0000010101000001: out_v[233] = 10'b0111101010;
    16'b1000010001000001: out_v[233] = 10'b0001111111;
    16'b0100110001000001: out_v[233] = 10'b1000110100;
    16'b0000010001000001: out_v[233] = 10'b0100011010;
    default: out_v[233] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1000000100000000: out_v[234] = 10'b1100001011;
    16'b1000000110000000: out_v[234] = 10'b0111001011;
    16'b1000001110000000: out_v[234] = 10'b0011100001;
    16'b1000000110000100: out_v[234] = 10'b0110001001;
    16'b1000000010000000: out_v[234] = 10'b1001001011;
    16'b0000001110000000: out_v[234] = 10'b1100110011;
    16'b0000001100000000: out_v[234] = 10'b0010011111;
    16'b1000000000000000: out_v[234] = 10'b1000110000;
    16'b0000000110000000: out_v[234] = 10'b1100100001;
    16'b1000001010000000: out_v[234] = 10'b0001011010;
    16'b0000000100000000: out_v[234] = 10'b0011101110;
    16'b1000001110000100: out_v[234] = 10'b0110100111;
    16'b0000001010000000: out_v[234] = 10'b1101000000;
    16'b1000000010000100: out_v[234] = 10'b0010011011;
    16'b0000000000000000: out_v[234] = 10'b0000111010;
    16'b1000001100000000: out_v[234] = 10'b0110100101;
    16'b1000001000000000: out_v[234] = 10'b0111000110;
    16'b0000000000000100: out_v[234] = 10'b0000000100;
    16'b0000001000000000: out_v[234] = 10'b0011001100;
    16'b0000001000000100: out_v[234] = 10'b0010101110;
    16'b0000000100000100: out_v[234] = 10'b0100001011;
    16'b0100000100000000: out_v[234] = 10'b0010001100;
    16'b0000000010000000: out_v[234] = 10'b0011110101;
    16'b0100000000000000: out_v[234] = 10'b1111001010;
    16'b1000000000000100: out_v[234] = 10'b0011011100;
    16'b0000001100000100: out_v[234] = 10'b0001001001;
    16'b1000000100000100: out_v[234] = 10'b1000110000;
    16'b0000010100000000: out_v[234] = 10'b0100111100;
    16'b0000000010010000: out_v[234] = 10'b0111010001;
    16'b0000000000010000: out_v[234] = 10'b1000111111;
    16'b1000000110000010: out_v[234] = 10'b1010000000;
    16'b1000011000000000: out_v[234] = 10'b1000011101;
    16'b1000001100000010: out_v[234] = 10'b1100100100;
    16'b1000000100000010: out_v[234] = 10'b1011000011;
    16'b1000001110000010: out_v[234] = 10'b1011011111;
    16'b0000001100000010: out_v[234] = 10'b1111111111;
    16'b1000001010010000: out_v[234] = 10'b1010001010;
    16'b0000001010010000: out_v[234] = 10'b1111100010;
    16'b0000001000010000: out_v[234] = 10'b1100000000;
    default: out_v[234] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000000101100: out_v[235] = 10'b0111001011;
    16'b0011000010001000: out_v[235] = 10'b0110100000;
    16'b0001000010001000: out_v[235] = 10'b0000011111;
    16'b0000000000101000: out_v[235] = 10'b0010100101;
    16'b0000000001101100: out_v[235] = 10'b1000111011;
    16'b0001000010000000: out_v[235] = 10'b1000010101;
    16'b0000000001001100: out_v[235] = 10'b1001011101;
    16'b0001000010101000: out_v[235] = 10'b1110111010;
    16'b0001000000001000: out_v[235] = 10'b0111010011;
    16'b0001000000101000: out_v[235] = 10'b0010011111;
    16'b0011000010101000: out_v[235] = 10'b1100100001;
    16'b0000000000100000: out_v[235] = 10'b1101100100;
    16'b0000000010101100: out_v[235] = 10'b0100011001;
    16'b0000000001100100: out_v[235] = 10'b1010011111;
    16'b0000000000100100: out_v[235] = 10'b1011000011;
    16'b0011000010000000: out_v[235] = 10'b1001100111;
    16'b0000000000001100: out_v[235] = 10'b0010111010;
    16'b0010000010101000: out_v[235] = 10'b0010011110;
    16'b0001000000101100: out_v[235] = 10'b0011011110;
    16'b0000000010101000: out_v[235] = 10'b0110001011;
    16'b0000000010001000: out_v[235] = 10'b1000011101;
    16'b0000000000001000: out_v[235] = 10'b1011111110;
    16'b0001000011101100: out_v[235] = 10'b1111011011;
    16'b0001000000000000: out_v[235] = 10'b1100011111;
    16'b0000000010100000: out_v[235] = 10'b1011001011;
    16'b0001000010101100: out_v[235] = 10'b0110010101;
    16'b0010000010001000: out_v[235] = 10'b0011100111;
    16'b0001000001101100: out_v[235] = 10'b1011110100;
    16'b0000000001101110: out_v[235] = 10'b1001110100;
    16'b0001000001001100: out_v[235] = 10'b0010111001;
    16'b0011000000001000: out_v[235] = 10'b0111100001;
    16'b0011000010100000: out_v[235] = 10'b1100110101;
    16'b0001000011001100: out_v[235] = 10'b1110111011;
    16'b0001000010100000: out_v[235] = 10'b0001011100;
    16'b0010000010100000: out_v[235] = 10'b0001101111;
    16'b0000000010001100: out_v[235] = 10'b1101100111;
    16'b0000000000001010: out_v[235] = 10'b0110111001;
    16'b0000000001001010: out_v[235] = 10'b1000100011;
    16'b0000000001000000: out_v[235] = 10'b0010011010;
    16'b0000000001000010: out_v[235] = 10'b0101000111;
    16'b0000000000000000: out_v[235] = 10'b1110100010;
    16'b0000000001001000: out_v[235] = 10'b0111011000;
    16'b0000000001101010: out_v[235] = 10'b1100000010;
    16'b0000000001000110: out_v[235] = 10'b0011010010;
    16'b0010000001000010: out_v[235] = 10'b0110010100;
    16'b0010000001000110: out_v[235] = 10'b0100000111;
    16'b0010000000001000: out_v[235] = 10'b0001011110;
    16'b0000000011101110: out_v[235] = 10'b1011000110;
    16'b0000000001001110: out_v[235] = 10'b1111000100;
    16'b0010000001100010: out_v[235] = 10'b0000011111;
    16'b0000000001100110: out_v[235] = 10'b0101110100;
    16'b0010000001100110: out_v[235] = 10'b0111000010;
    16'b0000000001101000: out_v[235] = 10'b0111010100;
    16'b0010000001000100: out_v[235] = 10'b1111110000;
    16'b0000000001100010: out_v[235] = 10'b0000111010;
    16'b0010000001001010: out_v[235] = 10'b1111000011;
    16'b0010000011101110: out_v[235] = 10'b0011111011;
    16'b0010000011001110: out_v[235] = 10'b0111101011;
    16'b0000000011001110: out_v[235] = 10'b0010101101;
    16'b0010000001101110: out_v[235] = 10'b0111011011;
    16'b0010000001001110: out_v[235] = 10'b1110010111;
    16'b0010000000101000: out_v[235] = 10'b1001001111;
    16'b0010000000000000: out_v[235] = 10'b1100011010;
    16'b0000000001100000: out_v[235] = 10'b0011111000;
    16'b0000000001000100: out_v[235] = 10'b1010101010;
    16'b0010000001100000: out_v[235] = 10'b0100001111;
    16'b0010000011001010: out_v[235] = 10'b0000101011;
    16'b0010000011100110: out_v[235] = 10'b0011011011;
    16'b0010000000001100: out_v[235] = 10'b0101011011;
    16'b0000000000000100: out_v[235] = 10'b0110101000;
    16'b0010000000000100: out_v[235] = 10'b0101011001;
    16'b0010000000101100: out_v[235] = 10'b0000011000;
    16'b0000000000001110: out_v[235] = 10'b1110111000;
    16'b0010000000100100: out_v[235] = 10'b0101011001;
    16'b0010000010000100: out_v[235] = 10'b1010010110;
    16'b0010000010001100: out_v[235] = 10'b1100110110;
    16'b0000000001100111: out_v[235] = 10'b0110100110;
    16'b0000000011100111: out_v[235] = 10'b0001101111;
    16'b0000000011000110: out_v[235] = 10'b1000001111;
    16'b0001000011100110: out_v[235] = 10'b0110010100;
    16'b0000000011100110: out_v[235] = 10'b1001010111;
    16'b1000000001100111: out_v[235] = 10'b0011011010;
    16'b0001000001101110: out_v[235] = 10'b0101111001;
    16'b0010000010101100: out_v[235] = 10'b0100100000;
    16'b0000000011100100: out_v[235] = 10'b1001001010;
    16'b0001000001100110: out_v[235] = 10'b0100010010;
    16'b0010000011000110: out_v[235] = 10'b0000001111;
    16'b0000000010100100: out_v[235] = 10'b1010011001;
    16'b0000000011101100: out_v[235] = 10'b0100110100;
    16'b1000000000001101: out_v[235] = 10'b0000110111;
    16'b0000000000001101: out_v[235] = 10'b0110011000;
    16'b0000000010000100: out_v[235] = 10'b1110011000;
    16'b0000000001001011: out_v[235] = 10'b1111011010;
    16'b1000000001001011: out_v[235] = 10'b1010001101;
    16'b0000000011001010: out_v[235] = 10'b1010101010;
    16'b0111000011100110: out_v[235] = 10'b1110110110;
    16'b0001000000100000: out_v[235] = 10'b1111001010;
    16'b0000000000100110: out_v[235] = 10'b1100110110;
    16'b0011000011100110: out_v[235] = 10'b1010001101;
    16'b0000000000101110: out_v[235] = 10'b0011110111;
    16'b0001000001100010: out_v[235] = 10'b1101001100;
    16'b0001000011100010: out_v[235] = 10'b1011101110;
    16'b0010001010000100: out_v[235] = 10'b1111010011;
    16'b0000000011000010: out_v[235] = 10'b0110111010;
    16'b0000000011000100: out_v[235] = 10'b1101111110;
    16'b0010000011000010: out_v[235] = 10'b0100011001;
    16'b0010000011000100: out_v[235] = 10'b0001110000;
    16'b0000000011101010: out_v[235] = 10'b0101011101;
    16'b0010000011101010: out_v[235] = 10'b1010011010;
    16'b0010000010100100: out_v[235] = 10'b0110101111;
    16'b0010001011100110: out_v[235] = 10'b0000110110;
    16'b0000000011001100: out_v[235] = 10'b1011001111;
    16'b0000001010100100: out_v[235] = 10'b0110100110;
    16'b0000001010000100: out_v[235] = 10'b1011000111;
    16'b0000001011100110: out_v[235] = 10'b1011100010;
    16'b0010001010100100: out_v[235] = 10'b0111110111;
    default: out_v[235] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1101100000100000: out_v[236] = 10'b1110011111;
    16'b1001100000001000: out_v[236] = 10'b0110001010;
    16'b1100100000100000: out_v[236] = 10'b1111000111;
    16'b1000100010101000: out_v[236] = 10'b0111010111;
    16'b0001100010100000: out_v[236] = 10'b0000111110;
    16'b0101100010100000: out_v[236] = 10'b0001011011;
    16'b0001100000000000: out_v[236] = 10'b1010111110;
    16'b1000100010100000: out_v[236] = 10'b1011010111;
    16'b1001101000001000: out_v[236] = 10'b0010010101;
    16'b0001100010000000: out_v[236] = 10'b1000000111;
    16'b0001100010100001: out_v[236] = 10'b0011011111;
    16'b1000100000100001: out_v[236] = 10'b1111010111;
    16'b1000000000100001: out_v[236] = 10'b1011010111;
    16'b1100100000100001: out_v[236] = 10'b1010010111;
    16'b1000100000101000: out_v[236] = 10'b1010000101;
    16'b0000100010000000: out_v[236] = 10'b1110000101;
    16'b1000000000100000: out_v[236] = 10'b0000111010;
    16'b0000100000100000: out_v[236] = 10'b1001010010;
    16'b0000100010100000: out_v[236] = 10'b1110011111;
    16'b1101100010100000: out_v[236] = 10'b0101100110;
    16'b1101100000100001: out_v[236] = 10'b1101010011;
    16'b0100100000100000: out_v[236] = 10'b1011010110;
    16'b0101100010100001: out_v[236] = 10'b0010000101;
    16'b1001101000101000: out_v[236] = 10'b0011110111;
    16'b0101100000100000: out_v[236] = 10'b0101111010;
    16'b1001100000000000: out_v[236] = 10'b1110011010;
    16'b0001100000100000: out_v[236] = 10'b1000001111;
    16'b1001100000101000: out_v[236] = 10'b1110000101;
    16'b0100100010100001: out_v[236] = 10'b0011010011;
    16'b0000100010001000: out_v[236] = 10'b0001010111;
    16'b0000000000100000: out_v[236] = 10'b0101100101;
    16'b1000100000100000: out_v[236] = 10'b1001010111;
    16'b1001100000100000: out_v[236] = 10'b1010111001;
    16'b1001100010101000: out_v[236] = 10'b1111101000;
    16'b0001100000001000: out_v[236] = 10'b1101110001;
    16'b1110100000100000: out_v[236] = 10'b1110010111;
    16'b0001100010101000: out_v[236] = 10'b1000111001;
    16'b1001001000001000: out_v[236] = 10'b0010011011;
    16'b1001100010100000: out_v[236] = 10'b1100100110;
    16'b1001100000100001: out_v[236] = 10'b0011000011;
    16'b0001100010001000: out_v[236] = 10'b0000011011;
    16'b0001100000101000: out_v[236] = 10'b1110011011;
    16'b1100100010100000: out_v[236] = 10'b0110001010;
    16'b1001000000100000: out_v[236] = 10'b1000011111;
    16'b0000100010101000: out_v[236] = 10'b0111111111;
    16'b1001000000000000: out_v[236] = 10'b1110001101;
    16'b0100100010100000: out_v[236] = 10'b1110011101;
    16'b1100000000100000: out_v[236] = 10'b0111011011;
    16'b0001001000000000: out_v[236] = 10'b1101000101;
    16'b0000001000000000: out_v[236] = 10'b1011001100;
    16'b0000000000000000: out_v[236] = 10'b0011000110;
    16'b0000000000001000: out_v[236] = 10'b1100100010;
    16'b0001000000000000: out_v[236] = 10'b0010100111;
    16'b0000001000001000: out_v[236] = 10'b0010110111;
    16'b0000001000000001: out_v[236] = 10'b0110111001;
    16'b0001001000000001: out_v[236] = 10'b0100110111;
    16'b0000000000001001: out_v[236] = 10'b1100111001;
    16'b0000001000001001: out_v[236] = 10'b1001001111;
    16'b1000001000000000: out_v[236] = 10'b1010010110;
    16'b0001001000001000: out_v[236] = 10'b0001110111;
    16'b0000000000000001: out_v[236] = 10'b1010001011;
    16'b1001001000000000: out_v[236] = 10'b1101010100;
    16'b1000000000000000: out_v[236] = 10'b0011000110;
    16'b0001000000000001: out_v[236] = 10'b1001110111;
    16'b0000001000101000: out_v[236] = 10'b0011001100;
    16'b0100001000001000: out_v[236] = 10'b1010010111;
    16'b1000101000001000: out_v[236] = 10'b0000011001;
    16'b0100001000000000: out_v[236] = 10'b1101101000;
    16'b0100000000000000: out_v[236] = 10'b0110000100;
    16'b0101000000000000: out_v[236] = 10'b0010011110;
    16'b1000101000000000: out_v[236] = 10'b1010010010;
    16'b0000101000100000: out_v[236] = 10'b1001110100;
    16'b1101101000101000: out_v[236] = 10'b0010010111;
    16'b1101001000101000: out_v[236] = 10'b1010110110;
    16'b0010001000001000: out_v[236] = 10'b1001010101;
    16'b0101101000001000: out_v[236] = 10'b1110111010;
    16'b1101101000001000: out_v[236] = 10'b0110001011;
    16'b1100101000001000: out_v[236] = 10'b0010100111;
    16'b0000001000100000: out_v[236] = 10'b1000100100;
    16'b0000101000101000: out_v[236] = 10'b1001101010;
    16'b1101101000000000: out_v[236] = 10'b0110101111;
    16'b0000101000001000: out_v[236] = 10'b0000010100;
    16'b1001001000101000: out_v[236] = 10'b1000100110;
    16'b0100001000101000: out_v[236] = 10'b0011000110;
    16'b1000001000001000: out_v[236] = 10'b0111111001;
    16'b0000101000000000: out_v[236] = 10'b0001000110;
    16'b0100101000001000: out_v[236] = 10'b0111001111;
    16'b1101001000001000: out_v[236] = 10'b0011101010;
    16'b1101001000100000: out_v[236] = 10'b1110011010;
    16'b1101001000000000: out_v[236] = 10'b1000011101;
    16'b1001101000000000: out_v[236] = 10'b0101011101;
    16'b0100000000001000: out_v[236] = 10'b1011010011;
    16'b0001101000001000: out_v[236] = 10'b0111110010;
    16'b0001001000101000: out_v[236] = 10'b0101110001;
    16'b0001101010001000: out_v[236] = 10'b1010111110;
    16'b1100001000001000: out_v[236] = 10'b0111111101;
    16'b0000100000001000: out_v[236] = 10'b0011100110;
    16'b0001101000000000: out_v[236] = 10'b0100110000;
    16'b0110000000000000: out_v[236] = 10'b1101000101;
    16'b1000101000101000: out_v[236] = 10'b1100010011;
    16'b0010001000101000: out_v[236] = 10'b1011110101;
    16'b0100001000000001: out_v[236] = 10'b1001011111;
    16'b0110001000000001: out_v[236] = 10'b1011010111;
    16'b1100001000000000: out_v[236] = 10'b1110101011;
    16'b0110001000110001: out_v[236] = 10'b0001010111;
    16'b0000001000100001: out_v[236] = 10'b0101110111;
    16'b0110001000010001: out_v[236] = 10'b1001010010;
    16'b0100001000100000: out_v[236] = 10'b1110100001;
    16'b0110000000010000: out_v[236] = 10'b0101011010;
    16'b0110001000110000: out_v[236] = 10'b0011011011;
    16'b0110001000100001: out_v[236] = 10'b0011001100;
    16'b0110000000010001: out_v[236] = 10'b0010001111;
    16'b1001001000000001: out_v[236] = 10'b1111001100;
    16'b1001001000100000: out_v[236] = 10'b0100001000;
    16'b0010001000000001: out_v[236] = 10'b1001110111;
    16'b0100000000000001: out_v[236] = 10'b1000011011;
    16'b1110001000000001: out_v[236] = 10'b1111000111;
    16'b0110001000000000: out_v[236] = 10'b0001101100;
    16'b0010000000000001: out_v[236] = 10'b0100100111;
    16'b0110001000010000: out_v[236] = 10'b1100011011;
    16'b0100001000100001: out_v[236] = 10'b1111110011;
    16'b1001000000001000: out_v[236] = 10'b1010111101;
    16'b0110000000000001: out_v[236] = 10'b0111110100;
    16'b0101001000000000: out_v[236] = 10'b0011111011;
    16'b1001001000100001: out_v[236] = 10'b0011011001;
    16'b1000001000100001: out_v[236] = 10'b0000110110;
    16'b0000000000100001: out_v[236] = 10'b0110011010;
    16'b0100000000100000: out_v[236] = 10'b0011111011;
    16'b0001001000100000: out_v[236] = 10'b0100111001;
    16'b1000101000001001: out_v[236] = 10'b0011011100;
    16'b1000001000101001: out_v[236] = 10'b1101011101;
    16'b0001101000100000: out_v[236] = 10'b1011001010;
    16'b0000001000101001: out_v[236] = 10'b1111000101;
    16'b1000101000100000: out_v[236] = 10'b0010111011;
    16'b0100101000100000: out_v[236] = 10'b1101111000;
    16'b1000001000101000: out_v[236] = 10'b1001001010;
    16'b0001101000101000: out_v[236] = 10'b1111011010;
    16'b1000001000001001: out_v[236] = 10'b1110000010;
    16'b1000101000101001: out_v[236] = 10'b1101011110;
    16'b1001101000100000: out_v[236] = 10'b1110000101;
    16'b1000001000100000: out_v[236] = 10'b0011011011;
    16'b1100101000100000: out_v[236] = 10'b1011001011;
    16'b0000101000101001: out_v[236] = 10'b1111100001;
    16'b1101101000100000: out_v[236] = 10'b0101011001;
    16'b0001001000101001: out_v[236] = 10'b0110111100;
    16'b0100000000100001: out_v[236] = 10'b0010110110;
    16'b1000001010001000: out_v[236] = 10'b0011100010;
    16'b0101001000100001: out_v[236] = 10'b0100010010;
    16'b1000101010001000: out_v[236] = 10'b1010101011;
    16'b0001000000101001: out_v[236] = 10'b0010011100;
    16'b0101000000100001: out_v[236] = 10'b0010100110;
    16'b0001000000100000: out_v[236] = 10'b0110110010;
    16'b0101001000100000: out_v[236] = 10'b1110100011;
    16'b0001001000100001: out_v[236] = 10'b0101111000;
    16'b0001000000100001: out_v[236] = 10'b0001100101;
    16'b0000000000101000: out_v[236] = 10'b1101101010;
    16'b0101000000100000: out_v[236] = 10'b0001110100;
    16'b1000000010000000: out_v[236] = 10'b1011111100;
    16'b0000000000101001: out_v[236] = 10'b0101011010;
    16'b1000000010001000: out_v[236] = 10'b0011110010;
    16'b0101101000101000: out_v[236] = 10'b0111010000;
    16'b0001000000001000: out_v[236] = 10'b1011101000;
    16'b0100101000101000: out_v[236] = 10'b1111100101;
    16'b0101101000100000: out_v[236] = 10'b1011010010;
    16'b0000100000101000: out_v[236] = 10'b0011111000;
    16'b1010001000111000: out_v[236] = 10'b0000100111;
    16'b1010001000101001: out_v[236] = 10'b0100111010;
    16'b1010000000110000: out_v[236] = 10'b1111010011;
    16'b1010001000110000: out_v[236] = 10'b1101101111;
    16'b1010001000111001: out_v[236] = 10'b0011111000;
    16'b1010001000101000: out_v[236] = 10'b0111000001;
    16'b0010001000111000: out_v[236] = 10'b1101000111;
    16'b1000001000111001: out_v[236] = 10'b0101110000;
    16'b0010001000110000: out_v[236] = 10'b1010101111;
    16'b1000001010101001: out_v[236] = 10'b1001111111;
    16'b1000000000110000: out_v[236] = 10'b1101111001;
    16'b0010001000101001: out_v[236] = 10'b1111100001;
    16'b0010001000100000: out_v[236] = 10'b0111100011;
    16'b0010001000111001: out_v[236] = 10'b1111111001;
    16'b1010000000110001: out_v[236] = 10'b0111010011;
    16'b1000001000111000: out_v[236] = 10'b0010111101;
    16'b1000001010101000: out_v[236] = 10'b0100110011;
    16'b1001000000101001: out_v[236] = 10'b1000011110;
    16'b1100001000100001: out_v[236] = 10'b1110110010;
    16'b1000000000101001: out_v[236] = 10'b0110100111;
    16'b1001001000101001: out_v[236] = 10'b0011011011;
    16'b0000001010100001: out_v[236] = 10'b0101000110;
    16'b1001001000001001: out_v[236] = 10'b1110101010;
    16'b0000001010101001: out_v[236] = 10'b0101011111;
    16'b1100001000100000: out_v[236] = 10'b1011010010;
    16'b0001001010101001: out_v[236] = 10'b0010011111;
    16'b1101001000100001: out_v[236] = 10'b1100011101;
    16'b0001001000001001: out_v[236] = 10'b0011010101;
    16'b1001001010101001: out_v[236] = 10'b1010110101;
    16'b1001000000000001: out_v[236] = 10'b0011111001;
    16'b1001000000001001: out_v[236] = 10'b1011110101;
    16'b1110001000100001: out_v[236] = 10'b1011111010;
    16'b1000101000100001: out_v[236] = 10'b1001100101;
    default: out_v[236] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010000011010100: out_v[237] = 10'b0100011011;
    16'b0010001010010100: out_v[237] = 10'b1011000011;
    16'b0001000000010100: out_v[237] = 10'b0110111011;
    16'b0010000000000100: out_v[237] = 10'b0011100010;
    16'b0010000010000100: out_v[237] = 10'b0110100011;
    16'b0000000010010100: out_v[237] = 10'b0001101000;
    16'b0000000011000100: out_v[237] = 10'b0101010011;
    16'b0000000000010100: out_v[237] = 10'b1100101110;
    16'b0010000010010100: out_v[237] = 10'b1100001001;
    16'b0011000010000100: out_v[237] = 10'b0101010111;
    16'b0000000010000100: out_v[237] = 10'b0011101001;
    16'b0000000000000100: out_v[237] = 10'b1110000101;
    16'b0010001010000100: out_v[237] = 10'b1011110010;
    16'b0010000000000000: out_v[237] = 10'b0010001111;
    16'b0010000011000100: out_v[237] = 10'b1000000011;
    16'b0001000000010000: out_v[237] = 10'b1001110011;
    16'b0011000000000100: out_v[237] = 10'b1111100100;
    16'b0011100000000000: out_v[237] = 10'b0000010001;
    16'b0001000000000000: out_v[237] = 10'b1010010001;
    16'b0001000000000100: out_v[237] = 10'b1111100110;
    16'b0010001011010100: out_v[237] = 10'b0001100111;
    16'b0011000000000000: out_v[237] = 10'b1001101001;
    16'b0000000011010100: out_v[237] = 10'b1101000001;
    16'b0010000001010000: out_v[237] = 10'b1000011111;
    16'b0001000010000100: out_v[237] = 10'b1111010011;
    16'b0011000010010100: out_v[237] = 10'b0110011110;
    16'b0011000000010100: out_v[237] = 10'b1001010111;
    16'b0010000000010100: out_v[237] = 10'b0111111011;
    16'b0000000000000000: out_v[237] = 10'b0001000101;
    16'b0001100000000000: out_v[237] = 10'b1100110101;
    16'b0000000001010000: out_v[237] = 10'b0111110011;
    16'b0010000011010000: out_v[237] = 10'b0011010001;
    16'b0010001100000000: out_v[237] = 10'b1011010111;
    16'b0010000100010000: out_v[237] = 10'b1100110101;
    16'b0000000100010000: out_v[237] = 10'b1100110111;
    16'b0000000100000000: out_v[237] = 10'b1010001100;
    16'b0010000100000000: out_v[237] = 10'b0011001111;
    16'b0000000110010100: out_v[237] = 10'b1010010010;
    16'b0000000000010000: out_v[237] = 10'b0010100111;
    16'b0010000101010000: out_v[237] = 10'b1101010010;
    16'b0010000000010000: out_v[237] = 10'b0101110100;
    16'b0000001100000000: out_v[237] = 10'b1100011111;
    16'b0010001100010000: out_v[237] = 10'b1100100111;
    16'b0000000100010100: out_v[237] = 10'b1000001110;
    16'b0000000101000000: out_v[237] = 10'b0011001100;
    16'b0010000101000000: out_v[237] = 10'b0010001011;
    16'b0001000100000000: out_v[237] = 10'b0101011110;
    16'b0000000001000000: out_v[237] = 10'b1100110100;
    16'b0001100100010000: out_v[237] = 10'b0000011010;
    16'b0010000001000000: out_v[237] = 10'b0111100110;
    16'b0010001101000000: out_v[237] = 10'b1001101010;
    16'b0000000100000100: out_v[237] = 10'b0111011110;
    16'b0001100100000000: out_v[237] = 10'b1011011010;
    16'b0001100001000000: out_v[237] = 10'b1101100100;
    16'b0000001001000000: out_v[237] = 10'b1110001101;
    16'b0001100101000000: out_v[237] = 10'b1001011010;
    16'b0001000101000000: out_v[237] = 10'b0001011011;
    16'b0001000001000000: out_v[237] = 10'b1011110000;
    16'b0011000100000000: out_v[237] = 10'b1001011100;
    16'b0011000001000000: out_v[237] = 10'b1101110110;
    16'b0011000101000000: out_v[237] = 10'b1110111001;
    16'b0010000101000100: out_v[237] = 10'b0001101100;
    16'b0000000101010000: out_v[237] = 10'b0111100000;
    16'b0010001001000000: out_v[237] = 10'b0001111010;
    16'b0011100101000000: out_v[237] = 10'b1000111100;
    16'b0010000001000100: out_v[237] = 10'b1000110011;
    16'b0001000100010000: out_v[237] = 10'b1011110001;
    16'b0000000110010000: out_v[237] = 10'b1101000111;
    16'b0100000100000000: out_v[237] = 10'b0011101000;
    16'b0000000011010000: out_v[237] = 10'b1100011011;
    16'b0010000111000000: out_v[237] = 10'b1010101111;
    16'b0000000111010100: out_v[237] = 10'b1101011001;
    16'b0000000111010000: out_v[237] = 10'b1000111100;
    16'b0001100101010000: out_v[237] = 10'b1000101111;
    16'b0001100111010100: out_v[237] = 10'b0110011011;
    16'b0010000111010100: out_v[237] = 10'b1111001100;
    16'b0000000111000000: out_v[237] = 10'b0110110110;
    16'b0010000111000100: out_v[237] = 10'b1101000110;
    16'b0010000111010000: out_v[237] = 10'b1001001100;
    16'b0000000111000100: out_v[237] = 10'b0100110010;
    16'b0001000101010000: out_v[237] = 10'b1011111100;
    16'b0000000001010100: out_v[237] = 10'b1100001101;
    16'b0000000101010100: out_v[237] = 10'b1010001111;
    16'b0100000111000100: out_v[237] = 10'b1001101011;
    16'b0010001111000100: out_v[237] = 10'b1100101100;
    16'b0000001111000100: out_v[237] = 10'b0011011011;
    16'b0000000101000100: out_v[237] = 10'b0110110111;
    16'b0010000110000100: out_v[237] = 10'b1001010101;
    16'b0000001011000100: out_v[237] = 10'b1110011110;
    16'b0001000111000100: out_v[237] = 10'b0100110110;
    16'b0000000110000100: out_v[237] = 10'b1111110000;
    16'b1000000111000100: out_v[237] = 10'b1111000000;
    16'b0011000111000100: out_v[237] = 10'b1101000001;
    16'b0110000111000100: out_v[237] = 10'b0001011111;
    16'b1001000101000000: out_v[237] = 10'b1010000001;
    16'b0000000001000100: out_v[237] = 10'b1001000010;
    16'b0000001101000100: out_v[237] = 10'b0011101110;
    16'b0000001111010100: out_v[237] = 10'b0100011010;
    16'b0000001001000100: out_v[237] = 10'b1101010100;
    16'b0100000011000100: out_v[237] = 10'b1111001110;
    16'b0011001111000100: out_v[237] = 10'b0111110001;
    16'b0010001011000100: out_v[237] = 10'b0101100011;
    16'b0010001110010100: out_v[237] = 10'b0010110111;
    16'b0010000110010100: out_v[237] = 10'b0011001101;
    16'b0010001110000100: out_v[237] = 10'b1101010101;
    16'b0100000010010100: out_v[237] = 10'b1001101111;
    16'b0010001111010100: out_v[237] = 10'b1011110000;
    16'b0000000010010000: out_v[237] = 10'b1110101100;
    16'b0010001000010000: out_v[237] = 10'b1001111001;
    16'b0001000101000100: out_v[237] = 10'b0111011110;
    16'b0001100011010100: out_v[237] = 10'b1101100101;
    16'b0100000001010100: out_v[237] = 10'b1100000111;
    16'b0001100001010100: out_v[237] = 10'b1010100011;
    16'b0100000011010100: out_v[237] = 10'b0111000100;
    16'b0101000001010100: out_v[237] = 10'b0000001110;
    16'b0101000011010100: out_v[237] = 10'b1001111110;
    16'b0001000001010100: out_v[237] = 10'b1010110111;
    16'b0101100001010000: out_v[237] = 10'b0111011011;
    16'b0100000111010100: out_v[237] = 10'b1001111111;
    16'b0101000101010000: out_v[237] = 10'b0000011011;
    16'b0101100101000000: out_v[237] = 10'b1111110000;
    16'b0101000001010000: out_v[237] = 10'b1101111011;
    16'b0001100101010100: out_v[237] = 10'b0011100110;
    16'b0100000101010000: out_v[237] = 10'b0111100001;
    16'b0101000100000000: out_v[237] = 10'b0000111100;
    16'b0100000101000000: out_v[237] = 10'b1111100010;
    16'b0101100001000000: out_v[237] = 10'b0110111010;
    16'b0001100001010000: out_v[237] = 10'b0011010111;
    16'b0100000001000000: out_v[237] = 10'b0100000010;
    16'b0100000001010000: out_v[237] = 10'b1111100101;
    16'b0101000001000000: out_v[237] = 10'b1100100111;
    16'b0101100001010100: out_v[237] = 10'b1001111001;
    16'b0100000100010000: out_v[237] = 10'b0010001000;
    16'b0101000101000000: out_v[237] = 10'b1101100011;
    16'b0001000001010000: out_v[237] = 10'b1010110101;
    16'b1001100001010100: out_v[237] = 10'b1100000110;
    16'b0101100101010100: out_v[237] = 10'b1011100110;
    16'b0101000101010100: out_v[237] = 10'b1111100111;
    16'b0101100100000000: out_v[237] = 10'b1011111010;
    16'b0001000101010100: out_v[237] = 10'b0110101111;
    16'b0101100101010000: out_v[237] = 10'b1101111011;
    16'b0001000011010100: out_v[237] = 10'b1000100011;
    16'b0101100011010100: out_v[237] = 10'b0011111111;
    16'b0001000110000100: out_v[237] = 10'b1010110111;
    16'b0010000100000100: out_v[237] = 10'b0111110011;
    16'b0010001101010000: out_v[237] = 10'b1111100010;
    16'b0001100111000100: out_v[237] = 10'b0101110010;
    16'b0000001110000100: out_v[237] = 10'b1101011001;
    16'b0010001100000100: out_v[237] = 10'b1111011011;
    16'b0010000101010100: out_v[237] = 10'b0111001010;
    16'b0010001101000100: out_v[237] = 10'b1111011100;
    16'b0011000110000100: out_v[237] = 10'b1010100011;
    16'b0100000101000100: out_v[237] = 10'b0000011111;
    16'b0100000110010100: out_v[237] = 10'b1011001001;
    16'b1000000111010100: out_v[237] = 10'b1001011111;
    16'b0110000111010100: out_v[237] = 10'b0011111100;
    16'b0100000110000100: out_v[237] = 10'b1001010001;
    16'b0110000101000100: out_v[237] = 10'b1101100101;
    16'b1001100101000000: out_v[237] = 10'b1001000111;
    16'b1001000001000000: out_v[237] = 10'b0101001010;
    16'b0100000001000100: out_v[237] = 10'b1101000111;
    16'b1001100001000000: out_v[237] = 10'b0111100011;
    default: out_v[237] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001000000000000: out_v[238] = 10'b0001011101;
    16'b0100101001000000: out_v[238] = 10'b1111101010;
    16'b1101101001000000: out_v[238] = 10'b1100111000;
    16'b0101101010000000: out_v[238] = 10'b1111010111;
    16'b0101100010000000: out_v[238] = 10'b0110011001;
    16'b0101101000000000: out_v[238] = 10'b1011000010;
    16'b1100101001000000: out_v[238] = 10'b0100101011;
    16'b1100001001000000: out_v[238] = 10'b1000011000;
    16'b0101001000000000: out_v[238] = 10'b1100100101;
    16'b1100101000000000: out_v[238] = 10'b0111111000;
    16'b0100101010000000: out_v[238] = 10'b1111101110;
    16'b0101101001000000: out_v[238] = 10'b0111011011;
    16'b0001101000000000: out_v[238] = 10'b1000100111;
    16'b0100101011000000: out_v[238] = 10'b0111110110;
    16'b0101101011000000: out_v[238] = 10'b0111101100;
    16'b1100100011000000: out_v[238] = 10'b0111011011;
    16'b1000001011000000: out_v[238] = 10'b1001010001;
    16'b1101101000000000: out_v[238] = 10'b1010111111;
    16'b1100101001000001: out_v[238] = 10'b0110000101;
    16'b0100100000000000: out_v[238] = 10'b1000010111;
    16'b0100100011000000: out_v[238] = 10'b1101101110;
    16'b0101100000000000: out_v[238] = 10'b0010011011;
    16'b0100100001000000: out_v[238] = 10'b1010011011;
    16'b0101000000000000: out_v[238] = 10'b0110000111;
    16'b1101101011000000: out_v[238] = 10'b0111101011;
    16'b1100100001000000: out_v[238] = 10'b0101001011;
    16'b0001001000000000: out_v[238] = 10'b0000011111;
    16'b1100101011000000: out_v[238] = 10'b0111000001;
    16'b1000101011000000: out_v[238] = 10'b0010111010;
    16'b0100001011000000: out_v[238] = 10'b1011110011;
    16'b1100001011000000: out_v[238] = 10'b1110001001;
    16'b0000000001000000: out_v[238] = 10'b1001111111;
    16'b0100100010000000: out_v[238] = 10'b1000111000;
    16'b0001100000000000: out_v[238] = 10'b1010010111;
    16'b1101101010000000: out_v[238] = 10'b1100110111;
    16'b0101001010000000: out_v[238] = 10'b1101011011;
    16'b0100101000000000: out_v[238] = 10'b1111001101;
    16'b1100101001100001: out_v[238] = 10'b1011000111;
    16'b0000001011000000: out_v[238] = 10'b1001000111;
    16'b0001000001000000: out_v[238] = 10'b1010110010;
    16'b0000000000100001: out_v[238] = 10'b1111010101;
    16'b1000000000100001: out_v[238] = 10'b0001100011;
    16'b1001000000100001: out_v[238] = 10'b1001110111;
    16'b0000000010100001: out_v[238] = 10'b1110010011;
    16'b1001000001100001: out_v[238] = 10'b0111000111;
    16'b1000000010100001: out_v[238] = 10'b1100010000;
    16'b0000001000100001: out_v[238] = 10'b0111000011;
    16'b1000000000100000: out_v[238] = 10'b1111000111;
    16'b1001000010100001: out_v[238] = 10'b1011001011;
    16'b1001000000100000: out_v[238] = 10'b1110010001;
    16'b0001000001100001: out_v[238] = 10'b1001011000;
    16'b1000000001100001: out_v[238] = 10'b1001001100;
    16'b0001000000100001: out_v[238] = 10'b0111000100;
    16'b0000001001000000: out_v[238] = 10'b0101000111;
    16'b1000001011100001: out_v[238] = 10'b0110101001;
    16'b1000001010100001: out_v[238] = 10'b0110101010;
    16'b1000001011100000: out_v[238] = 10'b1011011100;
    16'b0001001010100001: out_v[238] = 10'b0010110100;
    16'b1000001001000000: out_v[238] = 10'b0000110101;
    16'b0001000010100001: out_v[238] = 10'b1001000100;
    16'b1001001000100001: out_v[238] = 10'b1000101011;
    16'b1000000001000000: out_v[238] = 10'b1001000110;
    16'b1000100011000000: out_v[238] = 10'b1101101110;
    16'b1000101001000000: out_v[238] = 10'b1001110110;
    16'b1001001010100001: out_v[238] = 10'b1010110111;
    16'b1000001010000000: out_v[238] = 10'b0010010101;
    16'b1000001001100001: out_v[238] = 10'b1001100011;
    16'b1000001000100001: out_v[238] = 10'b0111110010;
    16'b1000000011010000: out_v[238] = 10'b0100111101;
    16'b0000000001100001: out_v[238] = 10'b0101011000;
    16'b1000000011000000: out_v[238] = 10'b1000001101;
    16'b1000100001000000: out_v[238] = 10'b1110001110;
    16'b1001001011000000: out_v[238] = 10'b1000111110;
    16'b1001000001000000: out_v[238] = 10'b1101000110;
    16'b1000001011000001: out_v[238] = 10'b1011000010;
    16'b0001001000100001: out_v[238] = 10'b1101010110;
    16'b0000001011100001: out_v[238] = 10'b1111100110;
    16'b1000001011010000: out_v[238] = 10'b0010010111;
    16'b1000001001000001: out_v[238] = 10'b0011110110;
    16'b1000000001000001: out_v[238] = 10'b1011110101;
    16'b0000001001100001: out_v[238] = 10'b0100010111;
    16'b1001000000000000: out_v[238] = 10'b0000101110;
    16'b1001000011000000: out_v[238] = 10'b1010110110;
    16'b0001000001100000: out_v[238] = 10'b1001110011;
    16'b0001000001100101: out_v[238] = 10'b0000011110;
    16'b0001001001100001: out_v[238] = 10'b0111011010;
    16'b1000000011100001: out_v[238] = 10'b1101111010;
    16'b0101000000100001: out_v[238] = 10'b1111100110;
    16'b0101100000100001: out_v[238] = 10'b1100100100;
    16'b0000000011100001: out_v[238] = 10'b0111100000;
    16'b0101000001100001: out_v[238] = 10'b1100100101;
    16'b0001100000100001: out_v[238] = 10'b0011001011;
    16'b0001000000100000: out_v[238] = 10'b1000111011;
    16'b0100000001100001: out_v[238] = 10'b0110011110;
    16'b0001100010100001: out_v[238] = 10'b1111011010;
    16'b0001000011100001: out_v[238] = 10'b0110001000;
    16'b0101101000100001: out_v[238] = 10'b1011001011;
    16'b0001001011100001: out_v[238] = 10'b0100001011;
    16'b0001101000100001: out_v[238] = 10'b1110000001;
    16'b0101000011100001: out_v[238] = 10'b1110100011;
    16'b1100000001100001: out_v[238] = 10'b1001011111;
    16'b0000000001100000: out_v[238] = 10'b0100101100;
    16'b0101000010100001: out_v[238] = 10'b1001011110;
    16'b1100000000000000: out_v[238] = 10'b1001111101;
    16'b0101000001000001: out_v[238] = 10'b0001011111;
    16'b1100000001100000: out_v[238] = 10'b1101010011;
    16'b1100100000100001: out_v[238] = 10'b0010111111;
    16'b0101000001100000: out_v[238] = 10'b0011110101;
    16'b0101000001000000: out_v[238] = 10'b0110101011;
    16'b1100000001000001: out_v[238] = 10'b0010011100;
    16'b0101100001100000: out_v[238] = 10'b0001110110;
    16'b1101000001100001: out_v[238] = 10'b1110001011;
    16'b0101100001000000: out_v[238] = 10'b0111001110;
    16'b1100000001000000: out_v[238] = 10'b1110101101;
    16'b0100000001000000: out_v[238] = 10'b1000011010;
    16'b0101100001100001: out_v[238] = 10'b0001010101;
    16'b0100100000100001: out_v[238] = 10'b1010011011;
    16'b1000000000000001: out_v[238] = 10'b0101110101;
    16'b1101000001000000: out_v[238] = 10'b1100010010;
    16'b0101000011000000: out_v[238] = 10'b0101001011;
    16'b0100100001100001: out_v[238] = 10'b1010101110;
    16'b0100000001100000: out_v[238] = 10'b1000101110;
    16'b1100000000100001: out_v[238] = 10'b1001010110;
    16'b1100100001100001: out_v[238] = 10'b0001110011;
    16'b1100100001100000: out_v[238] = 10'b1000111111;
    16'b1100100001000001: out_v[238] = 10'b1100011000;
    16'b0100000000000000: out_v[238] = 10'b0011110000;
    16'b1100000000000001: out_v[238] = 10'b0111100110;
    16'b1100100000000000: out_v[238] = 10'b0110010001;
    16'b1000000000000000: out_v[238] = 10'b0000111000;
    16'b0100000000100001: out_v[238] = 10'b0011111001;
    16'b0001000001000001: out_v[238] = 10'b0011111011;
    16'b1110000000000000: out_v[238] = 10'b0011011111;
    16'b0101100000000001: out_v[238] = 10'b0011110010;
    16'b1100001001100001: out_v[238] = 10'b0011101110;
    16'b0101000000100000: out_v[238] = 10'b1001100110;
    16'b1000001001100000: out_v[238] = 10'b0011011111;
    16'b0111000001000000: out_v[238] = 10'b1000100101;
    16'b0101001001100001: out_v[238] = 10'b1110000110;
    16'b1000000001100000: out_v[238] = 10'b1011111011;
    16'b0101100010100001: out_v[238] = 10'b1010101110;
    16'b1010000000000000: out_v[238] = 10'b1111011000;
    16'b1000001000100000: out_v[238] = 10'b1011011110;
    16'b1000000011110001: out_v[238] = 10'b0011001010;
    16'b1100101010110001: out_v[238] = 10'b0110111110;
    16'b0001000011010000: out_v[238] = 10'b0111011111;
    16'b1000000011110000: out_v[238] = 10'b1111100101;
    16'b1100101011100001: out_v[238] = 10'b0011100111;
    16'b0000000011010000: out_v[238] = 10'b0011101110;
    16'b1100101011010000: out_v[238] = 10'b0100001011;
    16'b1100100000100000: out_v[238] = 10'b0010101001;
    16'b1000100000100001: out_v[238] = 10'b1011101101;
    16'b1100101011110001: out_v[238] = 10'b0111000110;
    16'b1100101010010000: out_v[238] = 10'b1111110111;
    16'b0000000011110000: out_v[238] = 10'b0011111111;
    16'b1101100000100001: out_v[238] = 10'b0111101010;
    16'b1000100001100001: out_v[238] = 10'b0011101110;
    16'b0001000011000000: out_v[238] = 10'b1010100011;
    16'b0000000011110001: out_v[238] = 10'b1111011101;
    16'b1000001011110001: out_v[238] = 10'b1010011011;
    16'b1000100000000000: out_v[238] = 10'b0111101011;
    16'b1100101011110000: out_v[238] = 10'b1111001111;
    16'b1100101000100001: out_v[238] = 10'b1111101010;
    16'b1000101011010000: out_v[238] = 10'b1101000010;
    16'b1000000101000000: out_v[238] = 10'b0010001110;
    16'b1000000000000100: out_v[238] = 10'b0111100011;
    16'b1100010101000000: out_v[238] = 10'b1011011011;
    16'b0000010101000000: out_v[238] = 10'b1011100101;
    16'b1000000001000100: out_v[238] = 10'b0111100000;
    16'b1100000000000100: out_v[238] = 10'b0111001011;
    16'b1000010101000000: out_v[238] = 10'b0011101011;
    16'b1000000100000001: out_v[238] = 10'b0110011001;
    16'b1000000100000000: out_v[238] = 10'b0111110111;
    16'b1000100001000100: out_v[238] = 10'b1011100001;
    16'b1100000001000100: out_v[238] = 10'b0011110110;
    16'b0001010101000000: out_v[238] = 10'b1101011101;
    16'b1100000101000000: out_v[238] = 10'b0011111111;
    16'b0001010001000000: out_v[238] = 10'b1011110011;
    16'b0000000000100101: out_v[238] = 10'b1001000011;
    16'b1000000000100101: out_v[238] = 10'b1000001111;
    16'b1000010100000001: out_v[238] = 10'b0101110111;
    16'b1000010100100001: out_v[238] = 10'b1011100101;
    16'b1000010100000000: out_v[238] = 10'b1100100011;
    16'b0100010101000000: out_v[238] = 10'b0011001111;
    16'b0000000000000000: out_v[238] = 10'b0111001000;
    16'b1000010101100001: out_v[238] = 10'b0111100011;
    16'b1000010101000001: out_v[238] = 10'b1101110111;
    16'b0101010001000000: out_v[238] = 10'b0110101111;
    16'b0000000000000100: out_v[238] = 10'b0101011110;
    16'b1101000000100001: out_v[238] = 10'b0111010010;
    16'b1010001000100001: out_v[238] = 10'b0111001001;
    16'b1000001000000000: out_v[238] = 10'b1110110110;
    16'b1100000101100001: out_v[238] = 10'b1101010011;
    16'b1100010101100001: out_v[238] = 10'b1101011111;
    16'b1100000001100101: out_v[238] = 10'b1000000110;
    16'b0100010101100001: out_v[238] = 10'b1101100111;
    16'b0101010001100001: out_v[238] = 10'b0011100111;
    16'b1100000001100100: out_v[238] = 10'b1001111101;
    16'b1100000000100101: out_v[238] = 10'b1000111111;
    default: out_v[238] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1000011000000000: out_v[239] = 10'b0000011111;
    16'b1000011100000100: out_v[239] = 10'b0100010011;
    16'b1000011100100100: out_v[239] = 10'b0100111011;
    16'b1000010000000000: out_v[239] = 10'b1001101011;
    16'b1000010000100100: out_v[239] = 10'b0101001000;
    16'b1000010000000100: out_v[239] = 10'b1101000001;
    16'b0000010100000100: out_v[239] = 10'b1000011011;
    16'b1000000000000100: out_v[239] = 10'b0110011000;
    16'b0000010000000000: out_v[239] = 10'b0000100111;
    16'b1000011000000100: out_v[239] = 10'b0110010001;
    16'b1000010100000100: out_v[239] = 10'b1011000100;
    16'b1000001100000100: out_v[239] = 10'b0000010001;
    16'b1000010000000101: out_v[239] = 10'b1101000111;
    16'b0000010000000100: out_v[239] = 10'b1001110011;
    16'b1000011000000101: out_v[239] = 10'b0101100110;
    16'b0000010100100100: out_v[239] = 10'b1000110011;
    16'b0000010000000101: out_v[239] = 10'b0010101011;
    16'b0000011100100100: out_v[239] = 10'b1101111011;
    16'b1000110000000000: out_v[239] = 10'b0011011100;
    16'b0000011000100000: out_v[239] = 10'b1000101011;
    16'b1000010100100100: out_v[239] = 10'b1111001100;
    16'b1000111000000000: out_v[239] = 10'b0101010100;
    16'b0000011100000100: out_v[239] = 10'b0111110111;
    16'b1000001000000100: out_v[239] = 10'b0011100111;
    16'b1000011100000101: out_v[239] = 10'b1010011111;
    16'b1000111100100100: out_v[239] = 10'b0000011011;
    16'b0000011000000000: out_v[239] = 10'b1011000101;
    16'b1000011000100100: out_v[239] = 10'b1110000010;
    16'b1000111100000100: out_v[239] = 10'b1110111111;
    16'b0000011000000101: out_v[239] = 10'b1000111111;
    16'b0000111000000000: out_v[239] = 10'b1100010011;
    16'b0000000000000000: out_v[239] = 10'b1011000011;
    16'b0000100000000000: out_v[239] = 10'b0000011011;
    16'b0000110000100000: out_v[239] = 10'b1101001000;
    16'b0000110100000000: out_v[239] = 10'b1100001001;
    16'b0000110000000000: out_v[239] = 10'b1111001100;
    16'b0000100100000000: out_v[239] = 10'b0110010010;
    16'b0000111000100000: out_v[239] = 10'b1000001011;
    16'b0000110100100000: out_v[239] = 10'b1100010011;
    16'b0000010000100000: out_v[239] = 10'b1001000111;
    16'b0000110000000001: out_v[239] = 10'b1111010100;
    16'b1000110100000001: out_v[239] = 10'b0010101101;
    16'b0000110000000100: out_v[239] = 10'b1100011000;
    16'b0000010100100000: out_v[239] = 10'b0011011101;
    16'b1000110000100000: out_v[239] = 10'b0110110100;
    16'b0000010100000000: out_v[239] = 10'b0110110100;
    16'b1000110000000001: out_v[239] = 10'b0000111011;
    16'b1000110100000100: out_v[239] = 10'b1111001010;
    16'b1000110100100100: out_v[239] = 10'b1101010110;
    16'b0000100000000100: out_v[239] = 10'b0000110110;
    16'b1000010100100000: out_v[239] = 10'b1010100101;
    16'b0000011100000000: out_v[239] = 10'b0001011100;
    16'b1000110100100001: out_v[239] = 10'b1001010111;
    16'b1000010100100001: out_v[239] = 10'b0010100110;
    16'b0000110100000100: out_v[239] = 10'b1100011100;
    16'b1000100000100100: out_v[239] = 10'b1111110001;
    16'b1000100000100101: out_v[239] = 10'b0100110000;
    16'b1000110100000101: out_v[239] = 10'b0010101110;
    16'b1000010100000000: out_v[239] = 10'b1101011110;
    16'b1000100000000000: out_v[239] = 10'b0001101101;
    16'b1000100000000101: out_v[239] = 10'b1000110001;
    16'b0000011000000001: out_v[239] = 10'b1011011010;
    16'b1000100000000100: out_v[239] = 10'b1100110100;
    16'b1000110100100101: out_v[239] = 10'b1011010100;
    16'b0000010100000001: out_v[239] = 10'b0011010011;
    16'b1000110100000000: out_v[239] = 10'b1001111011;
    16'b1000010100000001: out_v[239] = 10'b1100110110;
    16'b1000010000000001: out_v[239] = 10'b1000111111;
    16'b1000000000000000: out_v[239] = 10'b0110011010;
    16'b1000110100100000: out_v[239] = 10'b0100110111;
    16'b1000111100100001: out_v[239] = 10'b1011110011;
    16'b0000010000000001: out_v[239] = 10'b0110101000;
    16'b1000110000100100: out_v[239] = 10'b0111011011;
    16'b1000111000000001: out_v[239] = 10'b0111000101;
    16'b1000110000000100: out_v[239] = 10'b0111101001;
    16'b0000110100100100: out_v[239] = 10'b1011100110;
    16'b1000100000000001: out_v[239] = 10'b0101010010;
    16'b0000111100000000: out_v[239] = 10'b0001101001;
    16'b1000011000000001: out_v[239] = 10'b1011010100;
    16'b1000110000100101: out_v[239] = 10'b0011011000;
    16'b1000110000000101: out_v[239] = 10'b0101001010;
    16'b1000001100000000: out_v[239] = 10'b0110011100;
    16'b1000011100000000: out_v[239] = 10'b0111101010;
    16'b1000101000000000: out_v[239] = 10'b1000110110;
    16'b1000101100000000: out_v[239] = 10'b0111010000;
    16'b1000001000000000: out_v[239] = 10'b0101111010;
    16'b1000111100100000: out_v[239] = 10'b0000011010;
    16'b1000011100000001: out_v[239] = 10'b0111011000;
    16'b0000111100100000: out_v[239] = 10'b0011110010;
    16'b1000111100000000: out_v[239] = 10'b0011111101;
    16'b1000111100000001: out_v[239] = 10'b1001110101;
    16'b1000011100100000: out_v[239] = 10'b0111011101;
    16'b0000001000000000: out_v[239] = 10'b1001101011;
    16'b0000001100000000: out_v[239] = 10'b1001100100;
    16'b0000101000000000: out_v[239] = 10'b0101010100;
    16'b0000011100100000: out_v[239] = 10'b1111011011;
    16'b0000101100000000: out_v[239] = 10'b0111010000;
    16'b1000101100000100: out_v[239] = 10'b0011001011;
    16'b0000111000000100: out_v[239] = 10'b1000110100;
    16'b0000000000000100: out_v[239] = 10'b1011010100;
    16'b1000000000000101: out_v[239] = 10'b1010111010;
    16'b0000100000100100: out_v[239] = 10'b1101101110;
    16'b0000101000000100: out_v[239] = 10'b1101101010;
    16'b0000011000000100: out_v[239] = 10'b0010011000;
    16'b1000101000000100: out_v[239] = 10'b1000111110;
    16'b1000010000100000: out_v[239] = 10'b0011110010;
    16'b0000111100000100: out_v[239] = 10'b1011111010;
    16'b1000111000000100: out_v[239] = 10'b1100111010;
    16'b1000011000100000: out_v[239] = 10'b0000111100;
    16'b1000111000100000: out_v[239] = 10'b0111001111;
    16'b0000110000100100: out_v[239] = 10'b0011000100;
    16'b0000010000100100: out_v[239] = 10'b0110100101;
    16'b0000000010000000: out_v[239] = 10'b1111101011;
    16'b0000000010010000: out_v[239] = 10'b0101000101;
    16'b0000000000010000: out_v[239] = 10'b1111111111;
    16'b0000001000000100: out_v[239] = 10'b0110111010;
    default: out_v[239] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001000001000000: out_v[240] = 10'b0110111010;
    16'b0100000001001000: out_v[240] = 10'b1100000001;
    16'b0001000001001000: out_v[240] = 10'b1110000000;
    16'b1101000001001000: out_v[240] = 10'b1010001101;
    16'b0000000000000000: out_v[240] = 10'b1001000100;
    16'b0001001000001000: out_v[240] = 10'b0100000111;
    16'b0001000000001000: out_v[240] = 10'b1001011000;
    16'b0000000000001000: out_v[240] = 10'b0101001000;
    16'b0101000001000000: out_v[240] = 10'b0101001010;
    16'b1001000001000000: out_v[240] = 10'b1100100110;
    16'b0000000001000000: out_v[240] = 10'b0001100011;
    16'b0101000000001000: out_v[240] = 10'b1100100011;
    16'b0101000001001000: out_v[240] = 10'b0100001001;
    16'b1001000001001000: out_v[240] = 10'b1010110010;
    16'b1000000001001000: out_v[240] = 10'b1000011011;
    16'b1001001000001000: out_v[240] = 10'b1011010001;
    16'b1001000000001000: out_v[240] = 10'b0001011010;
    16'b0000000001001000: out_v[240] = 10'b0100110110;
    16'b1101000001000000: out_v[240] = 10'b0101100000;
    16'b1001000000101000: out_v[240] = 10'b1000011111;
    16'b1001001001101000: out_v[240] = 10'b0100000110;
    16'b1101001001001000: out_v[240] = 10'b1100111111;
    16'b0100000001000000: out_v[240] = 10'b0101110111;
    16'b0100000000001000: out_v[240] = 10'b1100001101;
    16'b0001000000000000: out_v[240] = 10'b1010101100;
    16'b1001000000000000: out_v[240] = 10'b1111100010;
    16'b1001000001101000: out_v[240] = 10'b1111000000;
    16'b0101000000000000: out_v[240] = 10'b1100011010;
    16'b1001001000101000: out_v[240] = 10'b1011101011;
    16'b1101000000001000: out_v[240] = 10'b0110100011;
    16'b0100000000000000: out_v[240] = 10'b1000100110;
    16'b1001001001001000: out_v[240] = 10'b1100111010;
    16'b1000000001000000: out_v[240] = 10'b0011001100;
    16'b1000000000000000: out_v[240] = 10'b0010111010;
    16'b1000000000100000: out_v[240] = 10'b1000001110;
    16'b1000000001100000: out_v[240] = 10'b1011000101;
    16'b0001001000000000: out_v[240] = 10'b0001111110;
    16'b0000000000100000: out_v[240] = 10'b1100010100;
    16'b1100000000101000: out_v[240] = 10'b0010001111;
    16'b1100000000001000: out_v[240] = 10'b0010010100;
    16'b1000000000101000: out_v[240] = 10'b1110010010;
    16'b1001000000100000: out_v[240] = 10'b0101110011;
    16'b1000001000000000: out_v[240] = 10'b1110000111;
    16'b1000000000001000: out_v[240] = 10'b1110011011;
    16'b1001000001100000: out_v[240] = 10'b1001100100;
    16'b1100000000000000: out_v[240] = 10'b0010111100;
    16'b0000001000000000: out_v[240] = 10'b0011010110;
    16'b1000001001000000: out_v[240] = 10'b1011001111;
    16'b1001001000000000: out_v[240] = 10'b1001101100;
    16'b1100000001100000: out_v[240] = 10'b1011011111;
    16'b1100000001001000: out_v[240] = 10'b1000001001;
    16'b1100000000100000: out_v[240] = 10'b1101110001;
    16'b0100000000101000: out_v[240] = 10'b0111011100;
    16'b1100000001000000: out_v[240] = 10'b1110001010;
    16'b0100000000100000: out_v[240] = 10'b0110011100;
    16'b1000000001100001: out_v[240] = 10'b1011010010;
    16'b1000000000100001: out_v[240] = 10'b1100101001;
    16'b0001000000000001: out_v[240] = 10'b0011111111;
    16'b1001000000000001: out_v[240] = 10'b1000100111;
    16'b0001000000100000: out_v[240] = 10'b1111010011;
    16'b0000000000000001: out_v[240] = 10'b0001111010;
    16'b1101000000000000: out_v[240] = 10'b0101111001;
    16'b0001000000100001: out_v[240] = 10'b0111010011;
    16'b1101000001100000: out_v[240] = 10'b0001110100;
    16'b1001000001100001: out_v[240] = 10'b1000111101;
    16'b1101000001100001: out_v[240] = 10'b1010110111;
    16'b0001000000001001: out_v[240] = 10'b1110000000;
    16'b1001000000100001: out_v[240] = 10'b0100100000;
    16'b1000000000000001: out_v[240] = 10'b1001001111;
    16'b1001000000001001: out_v[240] = 10'b0000010010;
    default: out_v[240] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0111001001000000: out_v[241] = 10'b1011010101;
    16'b0111001000000000: out_v[241] = 10'b1101000110;
    16'b0101101001100000: out_v[241] = 10'b0010100010;
    16'b0110000000000000: out_v[241] = 10'b1001011110;
    16'b0001101000000000: out_v[241] = 10'b0011011111;
    16'b0010100000000000: out_v[241] = 10'b1110000011;
    16'b0101101001000000: out_v[241] = 10'b0110011110;
    16'b0000100000000000: out_v[241] = 10'b1000100101;
    16'b0101101001101000: out_v[241] = 10'b1100101011;
    16'b0001100000000000: out_v[241] = 10'b1110001011;
    16'b0111101001000000: out_v[241] = 10'b0001101111;
    16'b0111100000000000: out_v[241] = 10'b1001001111;
    16'b0111101001100000: out_v[241] = 10'b1010100001;
    16'b0110001001000000: out_v[241] = 10'b1001001111;
    16'b0111001001100000: out_v[241] = 10'b1110100110;
    16'b0011001001100000: out_v[241] = 10'b1010010111;
    16'b0001101000100000: out_v[241] = 10'b1100010111;
    16'b0001101001100000: out_v[241] = 10'b0101111001;
    16'b0100101001100000: out_v[241] = 10'b0110010111;
    16'b0011101001100000: out_v[241] = 10'b1001011110;
    16'b0101001001100000: out_v[241] = 10'b1011100010;
    16'b0110001001100000: out_v[241] = 10'b0100101111;
    16'b0110100000000000: out_v[241] = 10'b0001110100;
    16'b0111101001101000: out_v[241] = 10'b1101101011;
    16'b0111101000000000: out_v[241] = 10'b1101101101;
    16'b0011100000000000: out_v[241] = 10'b1110000111;
    16'b0110101001000000: out_v[241] = 10'b0011011011;
    16'b0101101000000000: out_v[241] = 10'b1110111110;
    16'b0010001001000000: out_v[241] = 10'b0000110011;
    16'b0010000000000000: out_v[241] = 10'b0000101101;
    16'b0110001000000000: out_v[241] = 10'b1101000100;
    16'b0111000000000000: out_v[241] = 10'b0101010110;
    16'b0110101000000000: out_v[241] = 10'b1110001010;
    16'b0001001001100000: out_v[241] = 10'b1100000111;
    16'b0011001001000000: out_v[241] = 10'b0001110110;
    16'b0101001001000000: out_v[241] = 10'b1011111110;
    16'b0101101000100000: out_v[241] = 10'b0101010110;
    16'b0001101001101000: out_v[241] = 10'b0111110001;
    16'b0100000000000000: out_v[241] = 10'b0101101011;
    16'b0000001000000000: out_v[241] = 10'b0100000110;
    16'b0000001001100000: out_v[241] = 10'b0110001001;
    16'b0000001001000000: out_v[241] = 10'b0000011111;
    16'b0000000000000000: out_v[241] = 10'b1011001000;
    16'b0000001000100000: out_v[241] = 10'b1000101000;
    16'b0000000000100000: out_v[241] = 10'b0010010110;
    16'b0100001000000000: out_v[241] = 10'b0110100101;
    16'b0100001001000000: out_v[241] = 10'b0110100100;
    16'b0001000000100000: out_v[241] = 10'b0001111011;
    16'b0001001001000000: out_v[241] = 10'b0101010011;
    16'b0001001001101000: out_v[241] = 10'b0110001100;
    16'b0101001001101000: out_v[241] = 10'b1100100010;
    16'b0100001001100000: out_v[241] = 10'b1001101100;
    16'b0010001001100000: out_v[241] = 10'b1101000101;
    16'b0100000001000000: out_v[241] = 10'b0100001000;
    16'b0000001001101000: out_v[241] = 10'b0101100101;
    16'b0100001001101000: out_v[241] = 10'b1000110100;
    16'b0101000001100000: out_v[241] = 10'b1111011011;
    16'b0101000000000000: out_v[241] = 10'b0010011110;
    16'b0001000000000000: out_v[241] = 10'b1100110100;
    16'b0101000001000000: out_v[241] = 10'b1110000110;
    16'b0101000001101000: out_v[241] = 10'b0101110110;
    16'b0011001001101000: out_v[241] = 10'b1010001111;
    16'b0100000001100000: out_v[241] = 10'b1011001101;
    16'b0101001000000000: out_v[241] = 10'b1001001100;
    16'b0111001001101000: out_v[241] = 10'b0010100110;
    16'b0001001011101000: out_v[241] = 10'b1101010110;
    16'b0001001001001000: out_v[241] = 10'b1101011111;
    16'b0001001000101000: out_v[241] = 10'b1000001101;
    16'b0000001000101000: out_v[241] = 10'b0111110000;
    16'b0011001000101000: out_v[241] = 10'b1101001001;
    16'b0010001001101000: out_v[241] = 10'b1110100001;
    16'b0010001011101000: out_v[241] = 10'b1100001010;
    16'b0110001001101000: out_v[241] = 10'b0111000010;
    16'b0111001011101000: out_v[241] = 10'b0011111001;
    16'b0010001000101000: out_v[241] = 10'b0111101110;
    16'b0001001000100000: out_v[241] = 10'b0101101110;
    16'b0011001011101000: out_v[241] = 10'b0001100110;
    16'b0011001000100000: out_v[241] = 10'b1001000010;
    16'b0010000000100000: out_v[241] = 10'b0001011010;
    16'b0010001000000000: out_v[241] = 10'b0011110110;
    16'b0111000000100000: out_v[241] = 10'b0110110011;
    16'b0001000000001000: out_v[241] = 10'b0011101110;
    16'b0000000000001000: out_v[241] = 10'b1110010000;
    16'b0110000000100000: out_v[241] = 10'b0000010000;
    16'b0010001000100000: out_v[241] = 10'b1010000100;
    16'b0011000000100000: out_v[241] = 10'b0001110001;
    16'b0011000000101000: out_v[241] = 10'b1110001011;
    16'b0101000000100000: out_v[241] = 10'b0101010110;
    16'b0011000000001000: out_v[241] = 10'b0011111011;
    16'b0010000000000001: out_v[241] = 10'b1110000000;
    16'b0011000000000000: out_v[241] = 10'b1110101001;
    16'b0101000000001000: out_v[241] = 10'b0011011011;
    16'b0010000000001000: out_v[241] = 10'b0011010011;
    16'b0111000000001000: out_v[241] = 10'b1110010101;
    16'b0111001000100000: out_v[241] = 10'b0111100110;
    16'b0011001000000000: out_v[241] = 10'b0111011010;
    16'b0110001000100000: out_v[241] = 10'b1111110011;
    16'b0011000001100000: out_v[241] = 10'b1001001110;
    16'b0001100000101000: out_v[241] = 10'b0000001100;
    16'b0011100000101000: out_v[241] = 10'b0111010000;
    16'b0010101001000000: out_v[241] = 10'b0001111010;
    16'b0011101001000000: out_v[241] = 10'b0011011100;
    16'b0001100000001000: out_v[241] = 10'b1111000010;
    16'b0001100001100000: out_v[241] = 10'b1111100110;
    16'b0011100000100000: out_v[241] = 10'b0111110010;
    16'b0001100000100000: out_v[241] = 10'b1111111011;
    16'b0000000000000001: out_v[241] = 10'b1010010011;
    16'b1001000100000000: out_v[241] = 10'b0100011100;
    16'b1001000000000000: out_v[241] = 10'b1110000000;
    16'b1000000000000000: out_v[241] = 10'b1011000010;
    16'b0001000100000000: out_v[241] = 10'b1111000011;
    16'b0100001000100001: out_v[241] = 10'b0011111011;
    16'b0100001000101000: out_v[241] = 10'b1011110111;
    16'b1011000000000000: out_v[241] = 10'b1010100010;
    16'b0100001000000001: out_v[241] = 10'b0000011101;
    16'b0000000000101000: out_v[241] = 10'b1111100001;
    16'b0100001000100000: out_v[241] = 10'b1011100011;
    16'b0000001000101001: out_v[241] = 10'b1110110010;
    16'b1010000000000000: out_v[241] = 10'b1010101111;
    16'b0000001000100001: out_v[241] = 10'b0110110011;
    16'b0110001000000001: out_v[241] = 10'b1001000011;
    16'b0110000000000001: out_v[241] = 10'b1011001110;
    16'b0001001000000000: out_v[241] = 10'b0000001111;
    16'b0011000100000000: out_v[241] = 10'b1101000111;
    16'b1011000100000000: out_v[241] = 10'b1101011111;
    default: out_v[241] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000100100001000: out_v[242] = 10'b0010010011;
    16'b0000000101001000: out_v[242] = 10'b1000110011;
    16'b0001100101001000: out_v[242] = 10'b1111111101;
    16'b0000100101001000: out_v[242] = 10'b1000110101;
    16'b0000000100101000: out_v[242] = 10'b0010111001;
    16'b0000100100001001: out_v[242] = 10'b1100001010;
    16'b0000000101101000: out_v[242] = 10'b0001100011;
    16'b0000100001000000: out_v[242] = 10'b0110110011;
    16'b0000100100101000: out_v[242] = 10'b1101110011;
    16'b0000000101001001: out_v[242] = 10'b0000010011;
    16'b0000100001001000: out_v[242] = 10'b1100010101;
    16'b0000100100101001: out_v[242] = 10'b0100111011;
    16'b0001100001001000: out_v[242] = 10'b0110000111;
    16'b0000000100001000: out_v[242] = 10'b0110010011;
    16'b0000100100000000: out_v[242] = 10'b0010100111;
    16'b0000000001001000: out_v[242] = 10'b1110001011;
    16'b0000100101000000: out_v[242] = 10'b1010100101;
    16'b0000100000000000: out_v[242] = 10'b0010110111;
    16'b0001100001000000: out_v[242] = 10'b1110001110;
    16'b0000000100000000: out_v[242] = 10'b1110011001;
    16'b0000000100101001: out_v[242] = 10'b1000000101;
    16'b0000100101001001: out_v[242] = 10'b0010001111;
    16'b0001000001001000: out_v[242] = 10'b0001001001;
    16'b0000000001000000: out_v[242] = 10'b1000011111;
    16'b0000100000001000: out_v[242] = 10'b0001101101;
    16'b0000000101101001: out_v[242] = 10'b0010000011;
    16'b0001100101001001: out_v[242] = 10'b1111011011;
    16'b0000000000101000: out_v[242] = 10'b1111001010;
    16'b0000000100001001: out_v[242] = 10'b1011101110;
    16'b0000000101000000: out_v[242] = 10'b0100100001;
    16'b0000000000001000: out_v[242] = 10'b0001101001;
    16'b0000100101101001: out_v[242] = 10'b0111101110;
    16'b0000100000001001: out_v[242] = 10'b0000100010;
    16'b0000100101000001: out_v[242] = 10'b0011110011;
    16'b0000000100100101: out_v[242] = 10'b0011010010;
    16'b0000000000000001: out_v[242] = 10'b1100101011;
    16'b0000000000000101: out_v[242] = 10'b1000101111;
    16'b0000000000100101: out_v[242] = 10'b0011110111;
    16'b0000000000100001: out_v[242] = 10'b1011000100;
    16'b0000000100000101: out_v[242] = 10'b0011100101;
    16'b0000100000101101: out_v[242] = 10'b0111000011;
    16'b0000000000101101: out_v[242] = 10'b0010011110;
    16'b0000000000001101: out_v[242] = 10'b0101010111;
    16'b0000000000000100: out_v[242] = 10'b1101000010;
    16'b0000100000101001: out_v[242] = 10'b1011010011;
    16'b0000000000000000: out_v[242] = 10'b1011110000;
    16'b0000000000101001: out_v[242] = 10'b1100011101;
    16'b0000100000100101: out_v[242] = 10'b0001111101;
    16'b0000000100100000: out_v[242] = 10'b1010000110;
    16'b0000100000100001: out_v[242] = 10'b1101001011;
    16'b0000000000100100: out_v[242] = 10'b1000101101;
    16'b0000100100000101: out_v[242] = 10'b1011100111;
    16'b0000000100100100: out_v[242] = 10'b0110110110;
    16'b0000100100100100: out_v[242] = 10'b1100001100;
    16'b0000100000000101: out_v[242] = 10'b0100000100;
    16'b0000000000100000: out_v[242] = 10'b0010100100;
    16'b0000100000100100: out_v[242] = 10'b1110110011;
    16'b0000000100000001: out_v[242] = 10'b0101011000;
    16'b0000100100100101: out_v[242] = 10'b1011001101;
    16'b0000100100100000: out_v[242] = 10'b0000110111;
    16'b0000100000100000: out_v[242] = 10'b1101100100;
    16'b0000100000000001: out_v[242] = 10'b0010111011;
    16'b0000100100000100: out_v[242] = 10'b1000010101;
    16'b0000000100000100: out_v[242] = 10'b0111001101;
    16'b0000100100101101: out_v[242] = 10'b0100111101;
    16'b0000100100000001: out_v[242] = 10'b1000011100;
    16'b0000100100101100: out_v[242] = 10'b1010010100;
    16'b0000000100101100: out_v[242] = 10'b1101000110;
    16'b0000000000101100: out_v[242] = 10'b0100100000;
    16'b0000100100100001: out_v[242] = 10'b1011001011;
    16'b0000000100100001: out_v[242] = 10'b1100001001;
    16'b0000000000001001: out_v[242] = 10'b0011111100;
    16'b0000100000101000: out_v[242] = 10'b0001010010;
    16'b0000000100101101: out_v[242] = 10'b1100010010;
    16'b0000100000101100: out_v[242] = 10'b1111101000;
    16'b0000101100100100: out_v[242] = 10'b0101000111;
    16'b0000101100100000: out_v[242] = 10'b1001101010;
    16'b0001000100101001: out_v[242] = 10'b0101100110;
    16'b0001000100101000: out_v[242] = 10'b0101101010;
    16'b0001000100101101: out_v[242] = 10'b0001100011;
    16'b0001000100001001: out_v[242] = 10'b1001111111;
    16'b0000000000001100: out_v[242] = 10'b0111101010;
    16'b0001000100100001: out_v[242] = 10'b1101110001;
    16'b0001000100001101: out_v[242] = 10'b1011000110;
    16'b0001000100101100: out_v[242] = 10'b0011010010;
    16'b0000000100001100: out_v[242] = 10'b0100010001;
    16'b0000100000000100: out_v[242] = 10'b1101001110;
    16'b0000100000001100: out_v[242] = 10'b0000110001;
    16'b0000100001100000: out_v[242] = 10'b1001011100;
    16'b0000100000001101: out_v[242] = 10'b0000001111;
    16'b0000000100101010: out_v[242] = 10'b0111000100;
    16'b0000000100100010: out_v[242] = 10'b1001100001;
    16'b0000010100100000: out_v[242] = 10'b0111100010;
    16'b0000000100101011: out_v[242] = 10'b0100001001;
    16'b0000010100101001: out_v[242] = 10'b1101001100;
    16'b0000000100100011: out_v[242] = 10'b1000101111;
    16'b0000010100101000: out_v[242] = 10'b0111110110;
    16'b0000010100100100: out_v[242] = 10'b0101001011;
    16'b0000010100100101: out_v[242] = 10'b0111100000;
    16'b0000000000100010: out_v[242] = 10'b0110110111;
    16'b0000010100101101: out_v[242] = 10'b0000101110;
    16'b0000010100101100: out_v[242] = 10'b0110001111;
    16'b0000000100101111: out_v[242] = 10'b0011001110;
    16'b0000000000100011: out_v[242] = 10'b0111111010;
    16'b0000000100001101: out_v[242] = 10'b0110010101;
    16'b0001000001101100: out_v[242] = 10'b0100011011;
    16'b0000100100001101: out_v[242] = 10'b0110011011;
    16'b0000000101101100: out_v[242] = 10'b1001001010;
    16'b0000101000100100: out_v[242] = 10'b0011101011;
    16'b0000000100101110: out_v[242] = 10'b1000101011;
    16'b0000101100101101: out_v[242] = 10'b1111000011;
    16'b0000000000101011: out_v[242] = 10'b1101100000;
    16'b0000101000100001: out_v[242] = 10'b1110000011;
    16'b0000101000100101: out_v[242] = 10'b1011111011;
    default: out_v[242] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010010001000010: out_v[243] = 10'b1000011100;
    16'b1000110000010000: out_v[243] = 10'b0011110011;
    16'b1110110101000010: out_v[243] = 10'b1000010001;
    16'b1010010101000010: out_v[243] = 10'b1001010110;
    16'b1000100000010000: out_v[243] = 10'b0010000111;
    16'b0110110101000010: out_v[243] = 10'b0011101110;
    16'b1100100000010000: out_v[243] = 10'b1011010111;
    16'b1010110101000010: out_v[243] = 10'b0010011011;
    16'b0001010001010010: out_v[243] = 10'b1110110001;
    16'b1110010101000010: out_v[243] = 10'b0011010111;
    16'b1110110101010010: out_v[243] = 10'b1000001111;
    16'b1000010001010010: out_v[243] = 10'b1001101110;
    16'b1100110101000010: out_v[243] = 10'b0111111010;
    16'b1000010001010000: out_v[243] = 10'b0011000100;
    16'b1100100100010000: out_v[243] = 10'b1100111011;
    16'b1110110101100010: out_v[243] = 10'b0000100101;
    16'b1001010000010000: out_v[243] = 10'b1100010101;
    16'b1000010000010000: out_v[243] = 10'b0101001111;
    16'b1100110101010010: out_v[243] = 10'b1010101110;
    16'b0110010101000010: out_v[243] = 10'b0010110100;
    16'b1110110001000010: out_v[243] = 10'b1010001111;
    16'b1100110101010000: out_v[243] = 10'b1101010101;
    16'b1100010101010010: out_v[243] = 10'b1101101001;
    16'b1000110001000010: out_v[243] = 10'b1010010111;
    16'b0001010001010000: out_v[243] = 10'b0011111101;
    16'b0010010101000010: out_v[243] = 10'b0100010110;
    16'b1010010001000010: out_v[243] = 10'b1010111001;
    16'b1110100101000010: out_v[243] = 10'b0010011111;
    16'b1000110001010010: out_v[243] = 10'b0111110101;
    16'b1110100101100010: out_v[243] = 10'b1010011111;
    16'b1100100101010000: out_v[243] = 10'b0001011010;
    16'b1100110001010000: out_v[243] = 10'b0011110101;
    16'b1010110001000010: out_v[243] = 10'b1011011010;
    16'b1000000000010000: out_v[243] = 10'b0100001010;
    16'b1110110100000010: out_v[243] = 10'b1000101010;
    16'b1000110001010000: out_v[243] = 10'b1111111110;
    16'b0001010000010000: out_v[243] = 10'b1000100110;
    16'b0000010001010010: out_v[243] = 10'b0001011001;
    16'b0000010001010000: out_v[243] = 10'b0011110001;
    16'b0000000000000000: out_v[243] = 10'b1100000111;
    16'b0000010000000000: out_v[243] = 10'b1100001011;
    16'b0000000001000000: out_v[243] = 10'b0011111000;
    16'b0000010001000000: out_v[243] = 10'b1110100001;
    16'b0000000001000010: out_v[243] = 10'b0110010111;
    16'b0000000001010010: out_v[243] = 10'b1011001000;
    16'b0010000001010010: out_v[243] = 10'b0101101101;
    16'b0000000001010000: out_v[243] = 10'b1000000111;
    16'b0000000000000010: out_v[243] = 10'b0000001110;
    16'b0010000001000010: out_v[243] = 10'b0000101100;
    16'b0001010000000000: out_v[243] = 10'b1001101001;
    16'b0000010000010000: out_v[243] = 10'b0111001100;
    16'b0001000000000000: out_v[243] = 10'b1001111101;
    16'b0000010001000010: out_v[243] = 10'b0101010110;
    16'b0010010001010010: out_v[243] = 10'b0000001010;
    16'b0001000001010000: out_v[243] = 10'b0101111101;
    16'b0011010001000010: out_v[243] = 10'b0001110001;
    16'b0000000001011000: out_v[243] = 10'b0010100010;
    16'b0001000001011000: out_v[243] = 10'b0111011011;
    16'b0000000101010000: out_v[243] = 10'b0111000111;
    16'b0001000000010000: out_v[243] = 10'b1101100001;
    16'b0001000101010000: out_v[243] = 10'b0101011110;
    16'b1000100001010000: out_v[243] = 10'b1011000010;
    16'b0011010101010010: out_v[243] = 10'b1111000101;
    16'b0000000000010000: out_v[243] = 10'b1001100100;
    16'b0001000101110000: out_v[243] = 10'b1100011111;
    16'b0001000001110000: out_v[243] = 10'b1100110001;
    16'b1001000001010000: out_v[243] = 10'b1111110011;
    16'b0001010101010000: out_v[243] = 10'b1000101100;
    16'b0010000000000010: out_v[243] = 10'b1110110101;
    16'b0001000001000000: out_v[243] = 10'b0010101100;
    16'b0000000101110000: out_v[243] = 10'b0111010111;
    16'b0001000000011000: out_v[243] = 10'b0110000110;
    16'b1001000101010000: out_v[243] = 10'b0011111011;
    16'b1000000001011000: out_v[243] = 10'b1010111011;
    16'b0011000001010010: out_v[243] = 10'b0010111110;
    16'b0011000001000010: out_v[243] = 10'b0001101000;
    16'b1000000001010000: out_v[243] = 10'b0011001111;
    16'b1001000001011000: out_v[243] = 10'b0000110111;
    16'b0000000100110000: out_v[243] = 10'b1100111100;
    16'b0011000101010010: out_v[243] = 10'b1011000011;
    16'b0011010001010010: out_v[243] = 10'b1010110110;
    16'b1011000001010010: out_v[243] = 10'b1001000110;
    16'b0000000001110000: out_v[243] = 10'b1110100100;
    16'b1001000000011000: out_v[243] = 10'b1010101111;
    16'b0011000001010000: out_v[243] = 10'b0111010101;
    16'b1001000000010000: out_v[243] = 10'b0011001111;
    16'b0011010101000010: out_v[243] = 10'b0010111010;
    16'b0010000101000010: out_v[243] = 10'b1101011111;
    16'b0111010001000010: out_v[243] = 10'b0110111011;
    16'b0010010101010010: out_v[243] = 10'b0001111000;
    16'b0001010101010010: out_v[243] = 10'b0001100110;
    16'b0000010101010010: out_v[243] = 10'b1100111010;
    16'b0001010001000010: out_v[243] = 10'b0101011100;
    16'b0010010000000010: out_v[243] = 10'b1110101011;
    16'b1011010001000010: out_v[243] = 10'b0001001010;
    16'b0011010000000010: out_v[243] = 10'b1001011001;
    16'b1001010001010000: out_v[243] = 10'b0110010011;
    16'b1011010101000010: out_v[243] = 10'b0000011101;
    16'b0111010101000010: out_v[243] = 10'b0101110110;
    16'b0110010001000010: out_v[243] = 10'b1010111011;
    16'b1011010101010010: out_v[243] = 10'b0111111010;
    16'b0111000100010010: out_v[243] = 10'b0011110001;
    16'b0111000100000000: out_v[243] = 10'b1101001111;
    16'b1101010101010000: out_v[243] = 10'b0001111101;
    16'b1101010000010000: out_v[243] = 10'b1101101001;
    16'b0111000100010000: out_v[243] = 10'b0111101101;
    16'b0001010001000000: out_v[243] = 10'b0110111001;
    16'b0111000000010010: out_v[243] = 10'b1010000000;
    16'b0001010100010000: out_v[243] = 10'b0111011011;
    16'b1101010100010000: out_v[243] = 10'b1010111010;
    16'b0001000001010010: out_v[243] = 10'b1000111001;
    16'b1111000100010010: out_v[243] = 10'b0010110011;
    16'b0011000100010010: out_v[243] = 10'b0111010010;
    16'b0101000100000000: out_v[243] = 10'b1101100011;
    16'b1001000000000000: out_v[243] = 10'b1001000111;
    16'b0101000100010000: out_v[243] = 10'b0101111101;
    16'b0011000100010000: out_v[243] = 10'b0011100011;
    16'b0011000000010010: out_v[243] = 10'b1000000100;
    16'b0101010000010000: out_v[243] = 10'b1100010111;
    16'b0101000100010010: out_v[243] = 10'b1001101111;
    16'b0101010100010000: out_v[243] = 10'b0010000110;
    16'b0001000100010000: out_v[243] = 10'b0011000011;
    16'b1101000000000000: out_v[243] = 10'b0011001100;
    16'b0001000000010010: out_v[243] = 10'b0110111001;
    16'b0001000100010010: out_v[243] = 10'b0011000100;
    16'b0101000000000000: out_v[243] = 10'b0101111011;
    16'b0111000101010010: out_v[243] = 10'b1111100010;
    16'b0101110100010000: out_v[243] = 10'b0111011111;
    16'b1101010100010010: out_v[243] = 10'b1111101001;
    16'b0111100100010010: out_v[243] = 10'b0110101101;
    16'b0010000100010010: out_v[243] = 10'b0011110000;
    16'b1101000100010010: out_v[243] = 10'b1000111111;
    16'b1000000000000000: out_v[243] = 10'b1100100000;
    16'b0010010000010010: out_v[243] = 10'b1111000000;
    16'b0000010000010010: out_v[243] = 10'b0111100100;
    16'b0110010100010010: out_v[243] = 10'b0110100111;
    16'b0110010100000010: out_v[243] = 10'b1001110111;
    16'b0111010101010010: out_v[243] = 10'b0001001101;
    16'b0010010100010010: out_v[243] = 10'b1000101001;
    16'b0100000000010000: out_v[243] = 10'b0110001100;
    16'b0110010101010010: out_v[243] = 10'b0101100100;
    16'b0111010100000010: out_v[243] = 10'b0100100011;
    16'b0011000101000010: out_v[243] = 10'b0001101111;
    16'b0010000001011010: out_v[243] = 10'b1011011011;
    16'b0001000001011010: out_v[243] = 10'b1110001100;
    16'b0010000001001010: out_v[243] = 10'b0011011101;
    16'b0001100101010000: out_v[243] = 10'b1100010111;
    16'b0000000000011000: out_v[243] = 10'b1011011001;
    16'b1101100100010000: out_v[243] = 10'b1111000110;
    16'b0101100101110000: out_v[243] = 10'b0011011011;
    16'b0001000000001010: out_v[243] = 10'b1001110011;
    16'b0001000000011010: out_v[243] = 10'b0110101011;
    16'b1001100101010000: out_v[243] = 10'b1110101010;
    16'b0000000000011010: out_v[243] = 10'b1110010110;
    16'b1101100101010000: out_v[243] = 10'b1011101011;
    16'b0001100001010000: out_v[243] = 10'b1010100111;
    16'b0001000000001000: out_v[243] = 10'b1011000101;
    16'b0101000101010000: out_v[243] = 10'b0000111001;
    16'b0001000001001010: out_v[243] = 10'b1001011000;
    16'b0000000000001000: out_v[243] = 10'b1110001010;
    16'b0001100000011000: out_v[243] = 10'b1111101000;
    16'b0000000001011010: out_v[243] = 10'b1011011111;
    16'b0101100101010000: out_v[243] = 10'b1100111100;
    16'b0010000000011010: out_v[243] = 10'b0011001000;
    16'b0001000001001000: out_v[243] = 10'b1101011011;
    16'b0011000001001010: out_v[243] = 10'b1110111111;
    16'b1001100001010000: out_v[243] = 10'b1001110100;
    16'b0001100001011000: out_v[243] = 10'b1110111111;
    16'b0000010100000000: out_v[243] = 10'b0011110000;
    16'b0101010100010010: out_v[243] = 10'b0011110111;
    16'b0000000100010000: out_v[243] = 10'b0001011100;
    16'b1001010100010000: out_v[243] = 10'b0110000111;
    16'b1000010100010000: out_v[243] = 10'b1011011011;
    16'b0000000100010010: out_v[243] = 10'b0010010001;
    16'b1001010100010010: out_v[243] = 10'b1101101111;
    16'b0000010100010000: out_v[243] = 10'b0000011111;
    16'b0001010100000000: out_v[243] = 10'b0011100001;
    16'b1001010101010000: out_v[243] = 10'b0011000100;
    16'b1001000100010000: out_v[243] = 10'b0001011101;
    16'b1001000100000000: out_v[243] = 10'b0011111111;
    16'b0001010100010010: out_v[243] = 10'b1101011011;
    16'b0001000100000000: out_v[243] = 10'b0011011111;
    16'b1110010101010010: out_v[243] = 10'b0011110111;
    16'b1000010101010010: out_v[243] = 10'b1010100111;
    16'b1011010001010010: out_v[243] = 10'b1001011001;
    16'b1010010001010010: out_v[243] = 10'b1110100111;
    16'b1010010101010010: out_v[243] = 10'b1001110110;
    16'b1001010000000000: out_v[243] = 10'b0110010000;
    16'b1111010101010010: out_v[243] = 10'b0111001011;
    16'b0000010101000000: out_v[243] = 10'b0111000001;
    16'b0110000101010010: out_v[243] = 10'b0110101110;
    16'b1001010001000000: out_v[243] = 10'b0101111110;
    16'b1111010101000010: out_v[243] = 10'b0101011001;
    16'b1000010000000000: out_v[243] = 10'b0111010111;
    16'b0000010101010000: out_v[243] = 10'b0110100000;
    16'b1001010101010010: out_v[243] = 10'b1011011111;
    16'b1001010001010010: out_v[243] = 10'b0111011101;
    16'b1000010001000000: out_v[243] = 10'b1111001011;
    16'b0010000101010010: out_v[243] = 10'b1100001011;
    16'b0101010101010010: out_v[243] = 10'b1010101000;
    16'b0101010101010000: out_v[243] = 10'b1011011110;
    16'b0111000101000000: out_v[243] = 10'b1111100010;
    16'b0001000101010010: out_v[243] = 10'b1011000010;
    16'b0111000101000010: out_v[243] = 10'b0110010010;
    16'b1111000101010010: out_v[243] = 10'b1010101111;
    16'b1101110100010000: out_v[243] = 10'b1000101011;
    16'b1101010101010010: out_v[243] = 10'b0100110010;
    16'b0101000101000000: out_v[243] = 10'b1011101111;
    16'b0101000101010010: out_v[243] = 10'b0011110111;
    16'b0000000000010010: out_v[243] = 10'b1101010111;
    16'b0111000101010000: out_v[243] = 10'b1000000111;
    default: out_v[243] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000000000000: out_v[244] = 10'b1010101001;
    16'b1000000000000001: out_v[244] = 10'b0000010001;
    16'b1000000000000000: out_v[244] = 10'b1001110001;
    16'b0000000000000001: out_v[244] = 10'b0111110001;
    16'b1000000010000000: out_v[244] = 10'b0000111101;
    16'b1000000000000101: out_v[244] = 10'b1111101100;
    16'b1000000000000100: out_v[244] = 10'b0101010100;
    16'b0000000000000100: out_v[244] = 10'b0100111010;
    16'b0000000010000100: out_v[244] = 10'b1111011010;
    16'b1000000010000100: out_v[244] = 10'b0111000000;
    16'b1100000000000100: out_v[244] = 10'b1001000110;
    16'b1100000000000000: out_v[244] = 10'b1111010111;
    16'b0100000000000100: out_v[244] = 10'b0101000101;
    16'b0000000010000000: out_v[244] = 10'b0010110111;
    16'b0000000010001100: out_v[244] = 10'b0010011000;
    16'b1010000000000100: out_v[244] = 10'b0010110111;
    16'b0010000000000000: out_v[244] = 10'b1000001010;
    16'b0000000010001000: out_v[244] = 10'b0110011011;
    16'b0010000000000100: out_v[244] = 10'b0001011011;
    16'b0000000000000101: out_v[244] = 10'b0100111000;
    16'b0000000100000100: out_v[244] = 10'b1101101011;
    16'b0000000000100000: out_v[244] = 10'b1010000011;
    16'b0000000010101000: out_v[244] = 10'b0111000101;
    16'b0000000010100000: out_v[244] = 10'b1100001101;
    default: out_v[244] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000110101000: out_v[245] = 10'b1110000001;
    16'b0000001101001011: out_v[245] = 10'b0011011111;
    16'b0000001101101011: out_v[245] = 10'b0001100110;
    16'b0000000111101010: out_v[245] = 10'b1100111100;
    16'b0000000110001010: out_v[245] = 10'b1101001111;
    16'b0000001001101011: out_v[245] = 10'b1011000101;
    16'b0000000110101010: out_v[245] = 10'b1010110001;
    16'b0100001111111011: out_v[245] = 10'b1010100111;
    16'b0000000111101011: out_v[245] = 10'b1110011011;
    16'b0000000100101011: out_v[245] = 10'b1101011011;
    16'b0100001001110011: out_v[245] = 10'b1111011111;
    16'b0000000101101011: out_v[245] = 10'b0010010111;
    16'b0100001101110011: out_v[245] = 10'b1111100110;
    16'b0000000100101010: out_v[245] = 10'b1000011101;
    16'b0000000100001010: out_v[245] = 10'b0001100111;
    16'b0000001001001011: out_v[245] = 10'b1001011010;
    16'b0100000111110010: out_v[245] = 10'b0110011111;
    16'b0000001000001011: out_v[245] = 10'b0010011111;
    16'b0100001101111011: out_v[245] = 10'b0111011111;
    16'b0000000101001011: out_v[245] = 10'b1010000111;
    16'b0000001011001011: out_v[245] = 10'b0110100011;
    16'b0000000101101010: out_v[245] = 10'b1011110110;
    16'b0100000111101010: out_v[245] = 10'b1110110111;
    16'b0100000101110011: out_v[245] = 10'b1011011001;
    16'b0100001111110011: out_v[245] = 10'b1010101011;
    16'b0000001111101011: out_v[245] = 10'b0111111010;
    16'b0000000100001011: out_v[245] = 10'b0000011010;
    16'b0100000110101010: out_v[245] = 10'b0010000011;
    16'b0000000010101010: out_v[245] = 10'b0011001011;
    16'b0100000111111010: out_v[245] = 10'b0101010110;
    16'b0000001111001011: out_v[245] = 10'b0000101111;
    16'b0000001011101011: out_v[245] = 10'b0110010001;
    16'b0100000101110010: out_v[245] = 10'b1001111011;
    16'b0000000110000000: out_v[245] = 10'b0011100011;
    16'b0000000110000010: out_v[245] = 10'b0110010101;
    16'b0000000000000010: out_v[245] = 10'b0110000111;
    16'b0000000000100010: out_v[245] = 10'b1001111011;
    16'b0000000000000000: out_v[245] = 10'b1111010100;
    16'b0000000010000000: out_v[245] = 10'b1010110110;
    16'b0000000000100000: out_v[245] = 10'b0011010101;
    16'b0000000010100010: out_v[245] = 10'b1100100110;
    16'b0100000000000010: out_v[245] = 10'b0010110101;
    16'b0100000000000000: out_v[245] = 10'b1101001011;
    16'b0100000000001010: out_v[245] = 10'b1001011011;
    16'b0000000010000010: out_v[245] = 10'b1011000001;
    16'b0000000000101010: out_v[245] = 10'b1010100111;
    16'b0000000010100000: out_v[245] = 10'b0100010011;
    16'b0100000000100010: out_v[245] = 10'b0010010001;
    16'b0100000000001000: out_v[245] = 10'b0001010011;
    16'b0000000110100010: out_v[245] = 10'b0101010100;
    16'b0100000010100010: out_v[245] = 10'b1100100011;
    16'b0100000101100011: out_v[245] = 10'b1010110111;
    16'b0100000110110010: out_v[245] = 10'b0010100100;
    16'b0000000110100000: out_v[245] = 10'b0010110101;
    16'b0100000000110010: out_v[245] = 10'b0001101000;
    16'b0100000110100010: out_v[245] = 10'b0010110010;
    16'b0100000010110010: out_v[245] = 10'b1000100111;
    16'b0000000111000001: out_v[245] = 10'b1111000110;
    16'b0100000110100011: out_v[245] = 10'b1011010111;
    16'b0000000110100001: out_v[245] = 10'b0001100110;
    16'b0100000010000010: out_v[245] = 10'b0100100100;
    16'b0100000110100000: out_v[245] = 10'b0011100100;
    16'b0100000100100011: out_v[245] = 10'b0111110100;
    16'b0000000110000001: out_v[245] = 10'b1110001101;
    16'b0100000100110010: out_v[245] = 10'b0100101100;
    16'b0100000010100000: out_v[245] = 10'b1110100111;
    16'b0100000110110011: out_v[245] = 10'b0000101001;
    16'b0100000110100001: out_v[245] = 10'b1110111011;
    16'b0100000010000000: out_v[245] = 10'b0110111101;
    16'b0100000111100011: out_v[245] = 10'b1110000110;
    16'b0000000110100011: out_v[245] = 10'b0000011010;
    16'b0100000111100010: out_v[245] = 10'b0010000011;
    16'b0000000100100011: out_v[245] = 10'b0010011011;
    16'b0100000110110001: out_v[245] = 10'b1111110011;
    16'b0000000100100001: out_v[245] = 10'b1011010110;
    16'b0100000100100010: out_v[245] = 10'b0011110000;
    16'b0000000100100010: out_v[245] = 10'b0011001001;
    16'b0100000010110000: out_v[245] = 10'b1111001110;
    16'b0100000110110000: out_v[245] = 10'b1111000110;
    16'b0000000010010000: out_v[245] = 10'b0100111011;
    16'b0000000111100001: out_v[245] = 10'b1001100001;
    16'b0000000110110010: out_v[245] = 10'b1010010101;
    16'b0100000000110000: out_v[245] = 10'b1011101010;
    16'b0100000000101000: out_v[245] = 10'b0001101110;
    16'b0100000101100010: out_v[245] = 10'b1111111110;
    16'b0100000000101010: out_v[245] = 10'b0011001110;
    16'b0100000000100000: out_v[245] = 10'b1010001001;
    16'b0100000001011010: out_v[245] = 10'b1000100111;
    16'b0100000000111010: out_v[245] = 10'b1111010001;
    16'b0000000100000010: out_v[245] = 10'b1001001010;
    16'b0100000100110000: out_v[245] = 10'b1010001000;
    16'b0100000001110010: out_v[245] = 10'b1000100111;
    16'b0100000101111010: out_v[245] = 10'b0101100000;
    16'b0100000100101010: out_v[245] = 10'b1010001111;
    16'b0100000001001010: out_v[245] = 10'b1100011101;
    16'b0100000100100000: out_v[245] = 10'b0101001011;
    16'b0100000001111010: out_v[245] = 10'b0010100011;
    16'b0100000001101010: out_v[245] = 10'b0110011011;
    16'b0100000000111000: out_v[245] = 10'b0111101101;
    16'b0100000000010000: out_v[245] = 10'b1001101101;
    16'b0100000100111010: out_v[245] = 10'b1001000101;
    16'b1000000000010000: out_v[245] = 10'b0011110111;
    16'b0000000101010010: out_v[245] = 10'b0111111011;
    16'b0100000101101010: out_v[245] = 10'b1000111110;
    16'b0100000010101010: out_v[245] = 10'b0110101000;
    16'b0000000100110010: out_v[245] = 10'b1000011111;
    16'b1000000100010000: out_v[245] = 10'b1000111110;
    16'b0000000100010010: out_v[245] = 10'b1101100011;
    16'b0000000000010000: out_v[245] = 10'b1010000101;
    16'b0000000000101000: out_v[245] = 10'b1111100001;
    16'b0000000101010000: out_v[245] = 10'b1011000001;
    16'b0000000100001000: out_v[245] = 10'b0101011111;
    16'b0000000100010000: out_v[245] = 10'b1011000010;
    16'b0000000000001010: out_v[245] = 10'b1000110100;
    16'b1000000100010010: out_v[245] = 10'b1100100011;
    16'b0000000000001000: out_v[245] = 10'b0110010101;
    16'b0100000100010000: out_v[245] = 10'b0101011111;
    16'b0000000010001000: out_v[245] = 10'b1101011010;
    16'b0100000100001000: out_v[245] = 10'b0000101100;
    16'b0000000100000000: out_v[245] = 10'b0101011010;
    16'b0000000000110000: out_v[245] = 10'b0011110010;
    16'b0000000111001010: out_v[245] = 10'b0101010110;
    16'b0000000110001000: out_v[245] = 10'b1010110101;
    16'b0000000111010000: out_v[245] = 10'b0010011010;
    16'b1000000100001010: out_v[245] = 10'b0111001101;
    16'b0100000100001010: out_v[245] = 10'b0111100100;
    16'b0000000111001001: out_v[245] = 10'b0101110010;
    16'b0000000110010000: out_v[245] = 10'b0101011000;
    16'b0000000101001010: out_v[245] = 10'b0100101001;
    16'b1000000100001000: out_v[245] = 10'b0011100111;
    16'b0000000010101000: out_v[245] = 10'b1110000001;
    16'b0100000110001000: out_v[245] = 10'b0000111010;
    16'b0000000010001010: out_v[245] = 10'b1001010100;
    16'b1000000000001010: out_v[245] = 10'b1001001101;
    16'b0000000100011000: out_v[245] = 10'b0111110111;
    16'b0000000110001011: out_v[245] = 10'b1011011010;
    16'b0000001100001010: out_v[245] = 10'b1001100110;
    16'b0000000000001011: out_v[245] = 10'b1111110011;
    16'b0000000010001011: out_v[245] = 10'b1111100100;
    16'b0100000011111010: out_v[245] = 10'b0010110010;
    16'b0000000000011010: out_v[245] = 10'b0110100010;
    16'b1000000000001000: out_v[245] = 10'b1010100100;
    16'b0000000000101011: out_v[245] = 10'b1010110010;
    16'b0000000001101010: out_v[245] = 10'b1111110001;
    16'b1000000000011000: out_v[245] = 10'b1001111111;
    16'b0000000001111010: out_v[245] = 10'b0000111110;
    16'b0000000011101010: out_v[245] = 10'b1101000011;
    16'b0100000011000010: out_v[245] = 10'b1000010101;
    16'b0100000011011010: out_v[245] = 10'b1001100001;
    16'b0100000010001010: out_v[245] = 10'b1010010000;
    16'b0100000011101010: out_v[245] = 10'b0000111010;
    16'b0100000111010010: out_v[245] = 10'b1011000111;
    16'b0000000011101011: out_v[245] = 10'b1101110010;
    16'b0100000011010000: out_v[245] = 10'b1111111011;
    16'b0100000011001010: out_v[245] = 10'b1100110111;
    16'b0000000011101000: out_v[245] = 10'b1010011011;
    16'b0100000011001000: out_v[245] = 10'b1000001001;
    16'b0000000011001011: out_v[245] = 10'b1011100010;
    16'b0000000011001010: out_v[245] = 10'b0000111001;
    16'b0100000011010010: out_v[245] = 10'b0101100110;
    16'b0100000011110010: out_v[245] = 10'b1001011000;
    16'b0100000111001010: out_v[245] = 10'b1111100010;
    16'b0000001100011010: out_v[245] = 10'b1010001111;
    16'b1000000100011010: out_v[245] = 10'b0110100110;
    16'b0000000100011010: out_v[245] = 10'b1010100110;
    16'b1000000100011000: out_v[245] = 10'b1100000000;
    16'b1000000000010010: out_v[245] = 10'b0010110101;
    16'b1000000100000010: out_v[245] = 10'b1111011011;
    16'b0000000110010010: out_v[245] = 10'b1111000010;
    16'b0000100100001000: out_v[245] = 10'b0111100110;
    16'b1000000000000010: out_v[245] = 10'b0110011010;
    16'b1000010100001100: out_v[245] = 10'b1101001010;
    16'b0000000000010010: out_v[245] = 10'b0010101101;
    16'b1000010100011100: out_v[245] = 10'b0101011110;
    16'b0100000110111000: out_v[245] = 10'b1111000011;
    16'b0000001110101010: out_v[245] = 10'b0011011100;
    16'b0000001110001010: out_v[245] = 10'b0100101110;
    16'b0000001010001010: out_v[245] = 10'b1100001010;
    16'b0100000110101000: out_v[245] = 10'b0111000011;
    16'b0100000110111010: out_v[245] = 10'b0111001111;
    16'b0000000110111000: out_v[245] = 10'b1111011011;
    16'b1000000110001000: out_v[245] = 10'b1101000110;
    16'b0000000110111010: out_v[245] = 10'b0001101111;
    16'b0000000100101000: out_v[245] = 10'b1100000011;
    16'b0100000010111010: out_v[245] = 10'b1111111000;
    16'b1000000110011000: out_v[245] = 10'b1101100110;
    16'b1000000110000000: out_v[245] = 10'b1001100111;
    16'b1000000100000000: out_v[245] = 10'b0001011110;
    16'b1000000110001010: out_v[245] = 10'b1101100110;
    16'b1000000000000000: out_v[245] = 10'b0101111101;
    default: out_v[245] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000010111001010: out_v[246] = 10'b0110101111;
    16'b0000010001101000: out_v[246] = 10'b1011001010;
    16'b0001010101101000: out_v[246] = 10'b0011101011;
    16'b0001010101001010: out_v[246] = 10'b0101011001;
    16'b0001010111001000: out_v[246] = 10'b0110100000;
    16'b0000010001001010: out_v[246] = 10'b0100001110;
    16'b0000010100001000: out_v[246] = 10'b1011011110;
    16'b0000010101001000: out_v[246] = 10'b0110110100;
    16'b0000000101001000: out_v[246] = 10'b0000110111;
    16'b0000010001001000: out_v[246] = 10'b1011101011;
    16'b0000010011001010: out_v[246] = 10'b0011101011;
    16'b0000010101101010: out_v[246] = 10'b1111110010;
    16'b0000010101000010: out_v[246] = 10'b0000010111;
    16'b0000010101001010: out_v[246] = 10'b1100100001;
    16'b0001010101101010: out_v[246] = 10'b1111000011;
    16'b0000010101000000: out_v[246] = 10'b0100010100;
    16'b0001010101001000: out_v[246] = 10'b0000100011;
    16'b0001010001000000: out_v[246] = 10'b0100001101;
    16'b0000010001000010: out_v[246] = 10'b1100011001;
    16'b0001010111001010: out_v[246] = 10'b0100010101;
    16'b0001010101000100: out_v[246] = 10'b1000101010;
    16'b0001000101001000: out_v[246] = 10'b1000100100;
    16'b0000010101101000: out_v[246] = 10'b0110100010;
    16'b0000010100100000: out_v[246] = 10'b1000101100;
    16'b0000010100101000: out_v[246] = 10'b0101001111;
    16'b0000010100101010: out_v[246] = 10'b1101110101;
    16'b0000010011000010: out_v[246] = 10'b1100010101;
    16'b0000010111001000: out_v[246] = 10'b0011110000;
    16'b0001010100100000: out_v[246] = 10'b1001110110;
    16'b0000010011001000: out_v[246] = 10'b1101000111;
    16'b0001010101000000: out_v[246] = 10'b0011110000;
    16'b0000010011000000: out_v[246] = 10'b1001000011;
    16'b0000010111101010: out_v[246] = 10'b1110001111;
    16'b0000010001000000: out_v[246] = 10'b0110111010;
    16'b0000010001100000: out_v[246] = 10'b1000100111;
    16'b0000000000000000: out_v[246] = 10'b0000100010;
    16'b0000000001000000: out_v[246] = 10'b0001111000;
    16'b0000010000000000: out_v[246] = 10'b0111010000;
    16'b0000010010000000: out_v[246] = 10'b1111000010;
    16'b0000000100000000: out_v[246] = 10'b1001000001;
    16'b0000010011100000: out_v[246] = 10'b1010101100;
    16'b0000000010000000: out_v[246] = 10'b0000100110;
    16'b0000010000100000: out_v[246] = 10'b0111111001;
    16'b0000000101000000: out_v[246] = 10'b1001100010;
    16'b0000010010000010: out_v[246] = 10'b1000000111;
    16'b0001010101000010: out_v[246] = 10'b0101010110;
    16'b0001010001000100: out_v[246] = 10'b1110010001;
    16'b0000010110001000: out_v[246] = 10'b1100110110;
    16'b0000010010001000: out_v[246] = 10'b0101110000;
    16'b0001010011001000: out_v[246] = 10'b0110010110;
    16'b0000000110001000: out_v[246] = 10'b0100010111;
    16'b0000010000000010: out_v[246] = 10'b1010000101;
    16'b0001010111001110: out_v[246] = 10'b0110010101;
    16'b0001010111000000: out_v[246] = 10'b1110010010;
    16'b0000010111000010: out_v[246] = 10'b1100000110;
    16'b0000010110001010: out_v[246] = 10'b1000000001;
    16'b0001010111000100: out_v[246] = 10'b1000111111;
    16'b0001000110001000: out_v[246] = 10'b1100100110;
    16'b0001010110001000: out_v[246] = 10'b1010010000;
    16'b0001010101001110: out_v[246] = 10'b0101000110;
    16'b0001010011000100: out_v[246] = 10'b1111011001;
    16'b0001010001001010: out_v[246] = 10'b1101010011;
    16'b0001010111000010: out_v[246] = 10'b0011100100;
    16'b0000010010001010: out_v[246] = 10'b0111110110;
    16'b0001010011000000: out_v[246] = 10'b1001010100;
    16'b0000010111000000: out_v[246] = 10'b0110011001;
    16'b0001010111001100: out_v[246] = 10'b1111010110;
    16'b0001010011001010: out_v[246] = 10'b1111110010;
    16'b0001010100101000: out_v[246] = 10'b0111010101;
    16'b0010010001001000: out_v[246] = 10'b0010110011;
    16'b0001010001001000: out_v[246] = 10'b1011001000;
    16'b0001010000101000: out_v[246] = 10'b1111000001;
    16'b0000010000101000: out_v[246] = 10'b0010001001;
    16'b0001010100001000: out_v[246] = 10'b1011101010;
    16'b0001010000100000: out_v[246] = 10'b1011011111;
    16'b0001000100001000: out_v[246] = 10'b1011001010;
    16'b0001010001101000: out_v[246] = 10'b1110010011;
    16'b0000010101100000: out_v[246] = 10'b0011101100;
    16'b0001010101100000: out_v[246] = 10'b0011011100;
    16'b0001010100101010: out_v[246] = 10'b1000111010;
    16'b0000000001001000: out_v[246] = 10'b1010001111;
    16'b0001010101001100: out_v[246] = 10'b1000110011;
    16'b0011010001001000: out_v[246] = 10'b1011110110;
    16'b0001010000001000: out_v[246] = 10'b0001001010;
    16'b0001000000101000: out_v[246] = 10'b1101100001;
    16'b0001000100000000: out_v[246] = 10'b1010001111;
    16'b0110010001001000: out_v[246] = 10'b0100110011;
    16'b0001010101100010: out_v[246] = 10'b1001110101;
    16'b0001000001001000: out_v[246] = 10'b0000101111;
    16'b0000000101100010: out_v[246] = 10'b0110011110;
    16'b0000010100000000: out_v[246] = 10'b1110100100;
    16'b0000000101000010: out_v[246] = 10'b0111111000;
    16'b0000000101100000: out_v[246] = 10'b0000111110;
    16'b0000000111100010: out_v[246] = 10'b0101111000;
    16'b0001000110000010: out_v[246] = 10'b1001111111;
    16'b0001000000000000: out_v[246] = 10'b1101101101;
    16'b0000000111000010: out_v[246] = 10'b0101111011;
    16'b0001010000000000: out_v[246] = 10'b0000111111;
    16'b0001000110001010: out_v[246] = 10'b0000111111;
    16'b0001010010001010: out_v[246] = 10'b0111110011;
    16'b0000000001100010: out_v[246] = 10'b0010111001;
    16'b0000000110000000: out_v[246] = 10'b0000111011;
    16'b0001000100000010: out_v[246] = 10'b0000110111;
    16'b0001000000001010: out_v[246] = 10'b1001001010;
    16'b0001010000001010: out_v[246] = 10'b1101000111;
    16'b0000000100000010: out_v[246] = 10'b0101011011;
    16'b0000000111001000: out_v[246] = 10'b1001011011;
    16'b0000000110001010: out_v[246] = 10'b0110010010;
    16'b0001010110000000: out_v[246] = 10'b0000111001;
    16'b0000010110000000: out_v[246] = 10'b1000111010;
    16'b0000000000001010: out_v[246] = 10'b0011100111;
    16'b0001000000000010: out_v[246] = 10'b1010111110;
    16'b0001010010001000: out_v[246] = 10'b0101011000;
    16'b0000000001000010: out_v[246] = 10'b1110000111;
    16'b0000000100001000: out_v[246] = 10'b1001100100;
    16'b0000000001100000: out_v[246] = 10'b0011010011;
    16'b0001010110001010: out_v[246] = 10'b1011000110;
    16'b0000000100001010: out_v[246] = 10'b0101001010;
    16'b0001000100001010: out_v[246] = 10'b0110110111;
    16'b0001000010001010: out_v[246] = 10'b0010111111;
    16'b0000000010001010: out_v[246] = 10'b1011101011;
    16'b0000000000000010: out_v[246] = 10'b0011011011;
    16'b0001010100000000: out_v[246] = 10'b0110110001;
    16'b0000010000001000: out_v[246] = 10'b0001110001;
    16'b0000000010000010: out_v[246] = 10'b1010010110;
    16'b0000000110000010: out_v[246] = 10'b1011001011;
    16'b0000000111001010: out_v[246] = 10'b0000100100;
    16'b0001010010000000: out_v[246] = 10'b0100011011;
    16'b0000000101001010: out_v[246] = 10'b1001101100;
    16'b0000000011000000: out_v[246] = 10'b1111101000;
    16'b0000010000001010: out_v[246] = 10'b0001111100;
    16'b0001000101000010: out_v[246] = 10'b1111001011;
    16'b0001010100001010: out_v[246] = 10'b1111100000;
    16'b0000100111001000: out_v[246] = 10'b1110011010;
    16'b0000100111001010: out_v[246] = 10'b1110010001;
    16'b0000000111000000: out_v[246] = 10'b1001011110;
    16'b0000000011001000: out_v[246] = 10'b1111000000;
    16'b0001000111001000: out_v[246] = 10'b1110000111;
    16'b0000100101001010: out_v[246] = 10'b1111110101;
    16'b0000100101001000: out_v[246] = 10'b1010101010;
    16'b0000100011001000: out_v[246] = 10'b1100011001;
    16'b0000100001001000: out_v[246] = 10'b1111000111;
    16'b0001000111000010: out_v[246] = 10'b0011010111;
    16'b0000100011001010: out_v[246] = 10'b1110110011;
    16'b0000110011001010: out_v[246] = 10'b1011011100;
    16'b0001001111001010: out_v[246] = 10'b1101001110;
    16'b0000110011001000: out_v[246] = 10'b0110010111;
    16'b0001000111001010: out_v[246] = 10'b1101001110;
    16'b0000000011001010: out_v[246] = 10'b1011101010;
    16'b0001000101001010: out_v[246] = 10'b0010100001;
    16'b0000010101100010: out_v[246] = 10'b1001001011;
    16'b0000010001100010: out_v[246] = 10'b1001100111;
    16'b0001010100000010: out_v[246] = 10'b1011110011;
    16'b0000010100001010: out_v[246] = 10'b1001000110;
    16'b0000010100000010: out_v[246] = 10'b1110100110;
    16'b0000000000001000: out_v[246] = 10'b0011001010;
    16'b0001000101100010: out_v[246] = 10'b0011111111;
    16'b0001000101000000: out_v[246] = 10'b1100010010;
    16'b0001000101100000: out_v[246] = 10'b0011101011;
    16'b0000010110100010: out_v[246] = 10'b0111101001;
    16'b0000010111100000: out_v[246] = 10'b1100000100;
    16'b0000010111100010: out_v[246] = 10'b1001100111;
    16'b0001010110100010: out_v[246] = 10'b1000101110;
    16'b0000010100100010: out_v[246] = 10'b0101110010;
    16'b0001010110100000: out_v[246] = 10'b0001101111;
    16'b0000010011100010: out_v[246] = 10'b1101111100;
    16'b0001010111100010: out_v[246] = 10'b0000110111;
    16'b0000010110100000: out_v[246] = 10'b0101010010;
    16'b0000000100100000: out_v[246] = 10'b1111000011;
    16'b0001010110101000: out_v[246] = 10'b0101110111;
    16'b0001010111101010: out_v[246] = 10'b0111011001;
    16'b0001010111100000: out_v[246] = 10'b1010011011;
    16'b0001010100100010: out_v[246] = 10'b0100111110;
    16'b0000010110000010: out_v[246] = 10'b1001000110;
    default: out_v[246] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000001100000: out_v[247] = 10'b1110000101;
    16'b0000100001101001: out_v[247] = 10'b0101000110;
    16'b0000100001101000: out_v[247] = 10'b1001000011;
    16'b0000010011000001: out_v[247] = 10'b1000000101;
    16'b0000000000100000: out_v[247] = 10'b1101001100;
    16'b0000110011101000: out_v[247] = 10'b1000111001;
    16'b0000100001001000: out_v[247] = 10'b0001110000;
    16'b0000000001000000: out_v[247] = 10'b1011100110;
    16'b0000000001101000: out_v[247] = 10'b1011100000;
    16'b0000100001001001: out_v[247] = 10'b0010110111;
    16'b0000100000001000: out_v[247] = 10'b1100100101;
    16'b0000000001001000: out_v[247] = 10'b1000100100;
    16'b0000010011000000: out_v[247] = 10'b0111011111;
    16'b0000000011100000: out_v[247] = 10'b1110001011;
    16'b0000000001000001: out_v[247] = 10'b0000001111;
    16'b0000000001001001: out_v[247] = 10'b0000101011;
    16'b0000000000000000: out_v[247] = 10'b1111000110;
    16'b0000110011001001: out_v[247] = 10'b1001000011;
    16'b0000100000001001: out_v[247] = 10'b0100101011;
    16'b0000110010001001: out_v[247] = 10'b1101000101;
    16'b0000000011000000: out_v[247] = 10'b0001011101;
    16'b0000100011101000: out_v[247] = 10'b0011011110;
    16'b0000000001100001: out_v[247] = 10'b0001110100;
    16'b0000010011001001: out_v[247] = 10'b1100011011;
    16'b0000110011101001: out_v[247] = 10'b1010111111;
    16'b0000010011100000: out_v[247] = 10'b0100011101;
    16'b0000100000101000: out_v[247] = 10'b0110010001;
    16'b0000000011101000: out_v[247] = 10'b0100101101;
    16'b0000100001100000: out_v[247] = 10'b1110011001;
    16'b1000000000000000: out_v[247] = 10'b0010100110;
    16'b0000010011101000: out_v[247] = 10'b0011000110;
    16'b1000000000100000: out_v[247] = 10'b0101011011;
    16'b1000000001100000: out_v[247] = 10'b1111000010;
    16'b0000000000100001: out_v[247] = 10'b1100000100;
    16'b0000000000000001: out_v[247] = 10'b1100001010;
    16'b0000010001100001: out_v[247] = 10'b0011110111;
    16'b0000010011100001: out_v[247] = 10'b1101001010;
    16'b0000110001101001: out_v[247] = 10'b1000111101;
    16'b0001000000000000: out_v[247] = 10'b1010101010;
    16'b1001000000000000: out_v[247] = 10'b0110011100;
    16'b1000000001000000: out_v[247] = 10'b0000111010;
    16'b0000010000000001: out_v[247] = 10'b1111111011;
    16'b0000110001001001: out_v[247] = 10'b0001001010;
    16'b0000010001000001: out_v[247] = 10'b0111001000;
    16'b0000010010000000: out_v[247] = 10'b1101101011;
    16'b0000000000001000: out_v[247] = 10'b0011011011;
    16'b0000100001000000: out_v[247] = 10'b0101011111;
    16'b0000100011001000: out_v[247] = 10'b0111010011;
    16'b0000100000000000: out_v[247] = 10'b0100100000;
    16'b0000100000000001: out_v[247] = 10'b1001111010;
    16'b0000100000100000: out_v[247] = 10'b1001100001;
    16'b0100100000100000: out_v[247] = 10'b0011001100;
    16'b0100000000100000: out_v[247] = 10'b1001100000;
    16'b0100000000000000: out_v[247] = 10'b0011100001;
    16'b0000000000100100: out_v[247] = 10'b0111001011;
    16'b0000000000010000: out_v[247] = 10'b1000001100;
    16'b1000000000010000: out_v[247] = 10'b1011111011;
    16'b0000001001001000: out_v[247] = 10'b0110010001;
    16'b1000000001001000: out_v[247] = 10'b1001000101;
    16'b0000000000101000: out_v[247] = 10'b0100010011;
    16'b0000000001101001: out_v[247] = 10'b0111110011;
    16'b0000100000101001: out_v[247] = 10'b1101011100;
    default: out_v[247] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001000000000011: out_v[248] = 10'b1101001001;
    16'b0001010010010011: out_v[248] = 10'b1000100000;
    16'b1001010010010011: out_v[248] = 10'b1010100000;
    16'b1100010010010001: out_v[248] = 10'b1011111111;
    16'b0000000010000011: out_v[248] = 10'b1111010100;
    16'b0001000010000011: out_v[248] = 10'b1100100011;
    16'b1101000010000011: out_v[248] = 10'b1010110001;
    16'b0001000010000010: out_v[248] = 10'b1100011001;
    16'b0101010010010011: out_v[248] = 10'b0011101110;
    16'b1001010000010011: out_v[248] = 10'b1000100111;
    16'b1101000000000001: out_v[248] = 10'b0110010101;
    16'b0001010010000011: out_v[248] = 10'b1001011011;
    16'b0000010010010011: out_v[248] = 10'b1110010001;
    16'b1101010010010011: out_v[248] = 10'b0000001111;
    16'b1100010010010011: out_v[248] = 10'b0110011111;
    16'b1101010010010001: out_v[248] = 10'b1011000010;
    16'b1001010010010001: out_v[248] = 10'b1110001001;
    16'b0001010000010011: out_v[248] = 10'b1101000100;
    16'b1101010000010011: out_v[248] = 10'b0110001011;
    16'b1001000000000001: out_v[248] = 10'b1010100001;
    16'b0000010010000011: out_v[248] = 10'b0100011011;
    16'b1000010010010011: out_v[248] = 10'b0011011101;
    16'b0001010010010010: out_v[248] = 10'b1010001111;
    16'b1001000010000011: out_v[248] = 10'b0101011011;
    16'b1100010000010001: out_v[248] = 10'b0100001110;
    16'b1001010010010010: out_v[248] = 10'b1001011111;
    16'b1000000000000001: out_v[248] = 10'b0100001001;
    16'b0000000000000011: out_v[248] = 10'b0100011001;
    16'b0000000010000010: out_v[248] = 10'b0011110010;
    16'b0001000000000010: out_v[248] = 10'b1000010101;
    16'b1001000010000001: out_v[248] = 10'b0100101110;
    16'b1101010000010001: out_v[248] = 10'b1110011110;
    16'b1000010010010001: out_v[248] = 10'b0000110110;
    16'b1001010010000011: out_v[248] = 10'b1010010110;
    16'b1100000000000001: out_v[248] = 10'b1110010011;
    16'b1101000000000011: out_v[248] = 10'b1101011110;
    16'b1101000000000000: out_v[248] = 10'b1100000101;
    16'b0001000000000000: out_v[248] = 10'b0010001010;
    16'b0000000000000000: out_v[248] = 10'b1000101101;
    16'b0001000010000000: out_v[248] = 10'b0001011011;
    16'b0000000010000000: out_v[248] = 10'b1011101001;
    16'b0000000000000001: out_v[248] = 10'b1111000101;
    16'b0001000000000001: out_v[248] = 10'b0000100111;
    16'b0001010000000001: out_v[248] = 10'b1011001001;
    16'b0000000000000010: out_v[248] = 10'b0011110110;
    16'b0000010000010001: out_v[248] = 10'b0101010110;
    16'b0000010000000001: out_v[248] = 10'b1111001101;
    16'b0001000010001000: out_v[248] = 10'b0100100100;
    16'b0001000000001000: out_v[248] = 10'b1011011100;
    16'b0101000010000000: out_v[248] = 10'b1110100010;
    16'b1101000010000010: out_v[248] = 10'b0010101110;
    16'b0000010010010001: out_v[248] = 10'b0011001111;
    16'b0101000000000000: out_v[248] = 10'b0110001111;
    16'b0101000010001000: out_v[248] = 10'b0010010101;
    16'b1000000010000001: out_v[248] = 10'b0101111111;
    16'b0000010010000001: out_v[248] = 10'b0100001100;
    16'b0000000010001001: out_v[248] = 10'b1010110110;
    16'b0001010010010001: out_v[248] = 10'b1010001000;
    16'b0101000010000001: out_v[248] = 10'b1101111001;
    16'b0001000010001001: out_v[248] = 10'b0110110110;
    16'b0000000010001000: out_v[248] = 10'b1011000101;
    16'b0100000000000001: out_v[248] = 10'b1110110001;
    16'b0100000000000000: out_v[248] = 10'b1000110101;
    16'b0000000010000001: out_v[248] = 10'b1000010111;
    16'b0001001010000000: out_v[248] = 10'b0101110101;
    16'b1101000010000000: out_v[248] = 10'b1101011100;
    16'b0101000010000010: out_v[248] = 10'b1000010110;
    16'b1001000010000000: out_v[248] = 10'b1000010110;
    16'b0001000010000001: out_v[248] = 10'b0011011010;
    16'b0100000010000001: out_v[248] = 10'b0011011110;
    16'b0001010000010001: out_v[248] = 10'b1111100101;
    16'b0100010010010001: out_v[248] = 10'b1001110111;
    16'b0101000010001001: out_v[248] = 10'b1111010110;
    16'b0101000000001000: out_v[248] = 10'b1010001111;
    16'b0100010010000001: out_v[248] = 10'b1110000111;
    16'b0001010010000001: out_v[248] = 10'b0111000011;
    16'b0000010110010001: out_v[248] = 10'b1011001011;
    16'b0100000010000000: out_v[248] = 10'b1101001100;
    16'b0000010010011001: out_v[248] = 10'b0001011110;
    16'b1001000000000000: out_v[248] = 10'b0100011111;
    16'b0101000000000010: out_v[248] = 10'b0111011100;
    16'b1001000010000010: out_v[248] = 10'b0110001001;
    16'b0100000000000010: out_v[248] = 10'b1001001110;
    16'b0001000010001010: out_v[248] = 10'b0111011000;
    16'b0001000000001010: out_v[248] = 10'b1110011110;
    16'b0101000000001010: out_v[248] = 10'b1100011111;
    16'b1000000010000000: out_v[248] = 10'b1111101011;
    16'b1001001010000000: out_v[248] = 10'b1001110110;
    16'b0000010000010011: out_v[248] = 10'b0000111001;
    16'b1000010000000001: out_v[248] = 10'b1001011011;
    16'b1000010000010001: out_v[248] = 10'b1000011011;
    16'b1000001000000000: out_v[248] = 10'b0111000101;
    16'b1000010010000001: out_v[248] = 10'b0111010101;
    16'b1001001000000000: out_v[248] = 10'b0011110001;
    16'b1000000010000011: out_v[248] = 10'b0110000101;
    16'b1000000000000000: out_v[248] = 10'b0000110010;
    16'b0000010000000011: out_v[248] = 10'b0110110000;
    16'b1000001000000001: out_v[248] = 10'b1101110101;
    16'b1000010010000011: out_v[248] = 10'b1010101100;
    16'b0000000000010001: out_v[248] = 10'b1011100101;
    16'b1000000010000010: out_v[248] = 10'b1110101100;
    16'b0001010000000010: out_v[248] = 10'b1001100110;
    16'b1001010010000010: out_v[248] = 10'b1000100111;
    16'b0001010010000010: out_v[248] = 10'b0001100110;
    16'b1101000000000010: out_v[248] = 10'b0110101011;
    16'b1000000000000010: out_v[248] = 10'b0010101100;
    16'b1100000000000000: out_v[248] = 10'b1011110010;
    16'b0001010000000011: out_v[248] = 10'b0111101100;
    16'b1001000000000010: out_v[248] = 10'b0111101110;
    16'b0000000000010011: out_v[248] = 10'b0110100011;
    16'b1100000000000010: out_v[248] = 10'b1111000111;
    16'b0000000010010011: out_v[248] = 10'b1011111010;
    16'b1001010000000010: out_v[248] = 10'b1100100111;
    16'b0100000010000010: out_v[248] = 10'b1101000110;
    16'b0001000110000010: out_v[248] = 10'b0001100110;
    16'b1100000010001000: out_v[248] = 10'b1011101011;
    16'b1100000010000000: out_v[248] = 10'b1011000010;
    16'b1100000010000010: out_v[248] = 10'b1000100111;
    16'b0000000110000010: out_v[248] = 10'b1000110001;
    16'b0001000110000000: out_v[248] = 10'b1011100000;
    16'b1000000010001000: out_v[248] = 10'b1110001011;
    16'b1001000000000011: out_v[248] = 10'b1011001001;
    16'b1001010000000011: out_v[248] = 10'b0011101111;
    16'b1011000010000011: out_v[248] = 10'b0101011111;
    16'b1011000010000010: out_v[248] = 10'b1011010010;
    16'b0001010000010010: out_v[248] = 10'b1111001110;
    16'b1001010010000001: out_v[248] = 10'b1100001001;
    16'b1001010000010001: out_v[248] = 10'b1100101110;
    default: out_v[248] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1010000000000001: out_v[249] = 10'b0111010000;
    16'b0011000000000110: out_v[249] = 10'b1000110011;
    16'b0011010000000110: out_v[249] = 10'b1110011111;
    16'b0111010000000010: out_v[249] = 10'b0110010011;
    16'b0010000000000100: out_v[249] = 10'b0100110111;
    16'b0111010000000110: out_v[249] = 10'b1010100111;
    16'b0001010000000010: out_v[249] = 10'b1101000110;
    16'b0001000000000110: out_v[249] = 10'b0110010111;
    16'b0001000000000010: out_v[249] = 10'b0111011011;
    16'b0011000000000000: out_v[249] = 10'b1110010011;
    16'b0011000000000010: out_v[249] = 10'b0101000010;
    16'b0010000000000000: out_v[249] = 10'b1010100100;
    16'b0011001000000000: out_v[249] = 10'b0000111011;
    16'b0010000000000010: out_v[249] = 10'b1001100111;
    16'b0010001000000010: out_v[249] = 10'b0110011001;
    16'b0011001000000010: out_v[249] = 10'b1011100011;
    16'b0011001000000110: out_v[249] = 10'b1111010011;
    16'b0001010000000110: out_v[249] = 10'b0100000110;
    16'b0001001000000000: out_v[249] = 10'b0111001110;
    16'b0001001000000010: out_v[249] = 10'b1100110001;
    16'b0000000000000100: out_v[249] = 10'b0110110011;
    16'b0010001000000000: out_v[249] = 10'b0011111001;
    16'b0011010000000010: out_v[249] = 10'b1101010011;
    16'b1001000000000111: out_v[249] = 10'b0111101111;
    16'b0011010000000100: out_v[249] = 10'b1000110011;
    16'b1011000000000111: out_v[249] = 10'b1000110011;
    16'b0101010100000010: out_v[249] = 10'b0110010111;
    16'b0011010000000000: out_v[249] = 10'b1101110111;
    16'b0000000000000000: out_v[249] = 10'b1010101001;
    16'b0010000000000110: out_v[249] = 10'b1001001000;
    16'b1010000000000011: out_v[249] = 10'b0010010100;
    16'b1011010000000111: out_v[249] = 10'b1110010001;
    16'b0101010000000010: out_v[249] = 10'b0000101100;
    16'b0011000000000100: out_v[249] = 10'b0011011001;
    16'b0000001000000000: out_v[249] = 10'b0010011001;
    16'b1000000000000101: out_v[249] = 10'b1011001001;
    16'b1010000000000101: out_v[249] = 10'b1100111001;
    16'b1010001000000101: out_v[249] = 10'b0011001000;
    16'b1111010000000111: out_v[249] = 10'b0100110001;
    16'b0001000000000000: out_v[249] = 10'b1011101010;
    16'b1000000000000001: out_v[249] = 10'b1111000011;
    16'b0001010000000000: out_v[249] = 10'b1110101101;
    16'b0101010000000110: out_v[249] = 10'b1111011000;
    16'b1010000000000111: out_v[249] = 10'b0101011100;
    16'b0000000000000010: out_v[249] = 10'b0000111011;
    16'b1010001000000001: out_v[249] = 10'b0111001011;
    16'b0001011000000010: out_v[249] = 10'b1110111101;
    16'b0000001000000100: out_v[249] = 10'b0001110010;
    16'b0000000000000101: out_v[249] = 10'b1000011101;
    16'b1000000000000011: out_v[249] = 10'b1010000111;
    16'b0000000000000001: out_v[249] = 10'b0011100010;
    16'b1000001000000101: out_v[249] = 10'b1001101100;
    16'b1000001000001101: out_v[249] = 10'b0010111101;
    16'b0001001000000100: out_v[249] = 10'b1100000111;
    16'b1000001000001001: out_v[249] = 10'b1111100100;
    16'b1000001000000001: out_v[249] = 10'b1100010101;
    16'b1001000000000101: out_v[249] = 10'b1010101101;
    16'b0001000000000100: out_v[249] = 10'b1111001110;
    16'b1001001000001101: out_v[249] = 10'b1110101010;
    16'b1001000000000001: out_v[249] = 10'b1001010101;
    16'b1001001000100101: out_v[249] = 10'b1111011110;
    16'b1101010000000111: out_v[249] = 10'b0011001100;
    16'b1000000000000111: out_v[249] = 10'b1100110001;
    16'b1101011000000111: out_v[249] = 10'b1110100110;
    16'b1101010000000101: out_v[249] = 10'b0110100011;
    16'b1001001000000101: out_v[249] = 10'b1110100110;
    16'b0001001000000101: out_v[249] = 10'b0111011101;
    16'b1001001000000111: out_v[249] = 10'b1110110100;
    16'b1000001000100101: out_v[249] = 10'b1101111100;
    16'b1001010000000101: out_v[249] = 10'b1110101100;
    16'b1000001000101101: out_v[249] = 10'b0110010110;
    16'b1000001000101001: out_v[249] = 10'b0001110011;
    16'b0000001000000101: out_v[249] = 10'b1011001110;
    16'b1001011000000101: out_v[249] = 10'b0110011101;
    16'b1000001000100001: out_v[249] = 10'b1111110110;
    16'b1000000000100101: out_v[249] = 10'b0010101100;
    16'b1001010000000001: out_v[249] = 10'b1101101110;
    16'b1101010000000011: out_v[249] = 10'b1010000110;
    16'b1001001000101101: out_v[249] = 10'b0100110110;
    16'b1101011000000101: out_v[249] = 10'b1110000110;
    16'b1001001000000001: out_v[249] = 10'b0001011100;
    16'b1101010000000001: out_v[249] = 10'b0101100111;
    16'b0010001000001000: out_v[249] = 10'b1010011010;
    16'b0000000010100000: out_v[249] = 10'b0010101010;
    16'b0010000010100000: out_v[249] = 10'b1010101101;
    16'b0000000010000000: out_v[249] = 10'b1010001011;
    16'b0010000000100000: out_v[249] = 10'b0000011101;
    16'b0000000000100000: out_v[249] = 10'b1101011111;
    16'b0010001000000100: out_v[249] = 10'b0100010111;
    16'b0010001000100000: out_v[249] = 10'b1011101011;
    16'b0101011000000000: out_v[249] = 10'b1110011010;
    16'b0010000010000000: out_v[249] = 10'b0011110100;
    16'b0000001000001000: out_v[249] = 10'b1010100011;
    16'b0010001000101000: out_v[249] = 10'b0110100101;
    16'b0000001000100000: out_v[249] = 10'b0010111011;
    16'b0000000000000110: out_v[249] = 10'b0010001001;
    16'b0000001000101000: out_v[249] = 10'b1011010001;
    16'b1010000010000001: out_v[249] = 10'b0110101110;
    16'b0010000000000111: out_v[249] = 10'b1010000100;
    16'b0010000000000101: out_v[249] = 10'b0100111000;
    16'b1011000000000101: out_v[249] = 10'b1101010011;
    16'b1011000000000001: out_v[249] = 10'b1101001010;
    16'b0010000000000001: out_v[249] = 10'b1010011110;
    16'b0101010000000100: out_v[249] = 10'b1110110110;
    16'b0001010000000100: out_v[249] = 10'b0001110111;
    16'b1011001000000101: out_v[249] = 10'b1011101010;
    16'b1011010000000101: out_v[249] = 10'b1011000010;
    16'b1010000000001101: out_v[249] = 10'b1011000010;
    16'b1010001000001101: out_v[249] = 10'b1010011011;
    16'b0000000000000111: out_v[249] = 10'b0111011001;
    16'b0000000100000000: out_v[249] = 10'b1011010110;
    16'b0000000000100100: out_v[249] = 10'b1011100111;
    16'b0000000010000100: out_v[249] = 10'b1100001101;
    16'b0000000100000110: out_v[249] = 10'b1110001100;
    16'b0000000110000000: out_v[249] = 10'b0110010101;
    16'b1001000000000011: out_v[249] = 10'b0010110101;
    16'b1000001000000011: out_v[249] = 10'b1010110011;
    16'b1000000010000011: out_v[249] = 10'b0111110111;
    16'b0010000010000100: out_v[249] = 10'b0111000101;
    16'b1000000010000001: out_v[249] = 10'b1100001101;
    16'b1010000010000011: out_v[249] = 10'b0110101010;
    16'b1000000010000101: out_v[249] = 10'b0000111111;
    16'b1010000010000101: out_v[249] = 10'b1000101011;
    default: out_v[249] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010100010010010: out_v[250] = 10'b1000001101;
    16'b0011100010000010: out_v[250] = 10'b0000011110;
    16'b0010100010000010: out_v[250] = 10'b1110001101;
    16'b0000100010010010: out_v[250] = 10'b1001110100;
    16'b0010000010010010: out_v[250] = 10'b1100110101;
    16'b0010100000010000: out_v[250] = 10'b1100000101;
    16'b0010000000010000: out_v[250] = 10'b1010001001;
    16'b0000110010000010: out_v[250] = 10'b1111110010;
    16'b0000100010000010: out_v[250] = 10'b0010100010;
    16'b0000000000010000: out_v[250] = 10'b1101001111;
    16'b0011100010010010: out_v[250] = 10'b0101000111;
    16'b0001100010000010: out_v[250] = 10'b0010110010;
    16'b0010100000010010: out_v[250] = 10'b0010010011;
    16'b0010110010000010: out_v[250] = 10'b0111100100;
    16'b0000000010010010: out_v[250] = 10'b0011001101;
    16'b0000100000000000: out_v[250] = 10'b1000110010;
    16'b0010100000000000: out_v[250] = 10'b1010001110;
    16'b0000110011000010: out_v[250] = 10'b0010011011;
    16'b0010110010010010: out_v[250] = 10'b1101101100;
    16'b0010110011000010: out_v[250] = 10'b1111101100;
    16'b0010100110010010: out_v[250] = 10'b0011001101;
    16'b0000100000010000: out_v[250] = 10'b1111000010;
    16'b0010100000000010: out_v[250] = 10'b1001011111;
    16'b0000000010000010: out_v[250] = 10'b0111011010;
    16'b0011110010000010: out_v[250] = 10'b0011110110;
    16'b0010000010000010: out_v[250] = 10'b0001111000;
    16'b0000000000000000: out_v[250] = 10'b1000011110;
    16'b0000000000000010: out_v[250] = 10'b1000101001;
    16'b0011100000010000: out_v[250] = 10'b0000110010;
    16'b0011000000010000: out_v[250] = 10'b0011111010;
    16'b0011100000000000: out_v[250] = 10'b1011001001;
    16'b0000100000000010: out_v[250] = 10'b1110111010;
    16'b0000000110010010: out_v[250] = 10'b1011010111;
    16'b0010000000000000: out_v[250] = 10'b0010111101;
    16'b0000100100010000: out_v[250] = 10'b1110000111;
    16'b0010101110010010: out_v[250] = 10'b0000110101;
    16'b0010100100010000: out_v[250] = 10'b1001011100;
    16'b0000000100010000: out_v[250] = 10'b1001110110;
    16'b0000100110010010: out_v[250] = 10'b0010100100;
    16'b0000100000010010: out_v[250] = 10'b1111100001;
    16'b0010100100000000: out_v[250] = 10'b0011111111;
    16'b0001000010000010: out_v[250] = 10'b1001001111;
    16'b0011100010000011: out_v[250] = 10'b0001011111;
    16'b0011000010000010: out_v[250] = 10'b1101100110;
    16'b0000000010000011: out_v[250] = 10'b1010011011;
    16'b0001100000000000: out_v[250] = 10'b1001101011;
    16'b0011100000000010: out_v[250] = 10'b1011001011;
    16'b0011000000000000: out_v[250] = 10'b0000011000;
    16'b0001000000000000: out_v[250] = 10'b0111011110;
    16'b0000000100000000: out_v[250] = 10'b1000010001;
    16'b0001000000010000: out_v[250] = 10'b0010110011;
    16'b0010000000000010: out_v[250] = 10'b0001111010;
    16'b0000010001000000: out_v[250] = 10'b0000101101;
    16'b0000010001010000: out_v[250] = 10'b1001101111;
    16'b0000010000010000: out_v[250] = 10'b0101101010;
    16'b0000100100000000: out_v[250] = 10'b0111100011;
    16'b0010010001010000: out_v[250] = 10'b1110010100;
    16'b0010010011000010: out_v[250] = 10'b0011110110;
    16'b1000000010010010: out_v[250] = 10'b1111011010;
    16'b0000000000010010: out_v[250] = 10'b1111010010;
    16'b0010000010000011: out_v[250] = 10'b0111100100;
    16'b0010000000000100: out_v[250] = 10'b1000001110;
    16'b0000000000000001: out_v[250] = 10'b0011010011;
    16'b0010000000000001: out_v[250] = 10'b1001110100;
    16'b0011000000000001: out_v[250] = 10'b1000111011;
    16'b0010000010000110: out_v[250] = 10'b1001111101;
    16'b0010000010000111: out_v[250] = 10'b1100010001;
    16'b0001100000010000: out_v[250] = 10'b1101000000;
    16'b0001100010010010: out_v[250] = 10'b1100000010;
    16'b0011110011010010: out_v[250] = 10'b1111010001;
    default: out_v[250] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000100000000000: out_v[251] = 10'b0101110010;
    16'b0000100001010000: out_v[251] = 10'b0010010011;
    16'b0000001011010001: out_v[251] = 10'b0011110100;
    16'b0000000000010000: out_v[251] = 10'b1000100110;
    16'b0000000000010100: out_v[251] = 10'b1011000110;
    16'b0000100010010001: out_v[251] = 10'b1100111010;
    16'b0000000001001001: out_v[251] = 10'b1100111011;
    16'b0000000000001000: out_v[251] = 10'b0111100011;
    16'b0000000000101100: out_v[251] = 10'b0111000011;
    16'b0000100001010001: out_v[251] = 10'b1101001101;
    16'b0000101011010001: out_v[251] = 10'b0100101110;
    16'b0000100000010000: out_v[251] = 10'b0111110011;
    16'b0000000000000000: out_v[251] = 10'b0110000111;
    16'b0000000000110000: out_v[251] = 10'b1111110011;
    16'b0000000001010000: out_v[251] = 10'b1110001111;
    16'b0000000000010001: out_v[251] = 10'b1110011111;
    16'b0000100001000000: out_v[251] = 10'b0101110010;
    16'b0000000000010101: out_v[251] = 10'b0110001011;
    16'b0000000000001001: out_v[251] = 10'b0111101100;
    16'b0000000000110100: out_v[251] = 10'b1110010101;
    16'b0000000000011000: out_v[251] = 10'b0110111110;
    16'b0000000011010001: out_v[251] = 10'b1011000011;
    16'b0000000001010001: out_v[251] = 10'b0100001111;
    16'b0000000000111100: out_v[251] = 10'b1101000011;
    16'b0000100000011001: out_v[251] = 10'b0000100110;
    16'b0000100000001001: out_v[251] = 10'b1110000111;
    16'b0000100001000001: out_v[251] = 10'b1110111110;
    16'b0000000000001100: out_v[251] = 10'b0001011011;
    16'b0000101010010001: out_v[251] = 10'b0111010001;
    16'b0000000010010001: out_v[251] = 10'b1001111110;
    16'b0000000001000000: out_v[251] = 10'b1100101110;
    16'b0000100011010001: out_v[251] = 10'b1001101011;
    16'b0000100000010001: out_v[251] = 10'b0111011001;
    16'b0000001010010001: out_v[251] = 10'b1101111001;
    16'b0000100001011001: out_v[251] = 10'b0111100010;
    16'b0000000000011001: out_v[251] = 10'b1011111110;
    16'b0000000000100000: out_v[251] = 10'b1010100100;
    16'b0000000000100100: out_v[251] = 10'b1001100010;
    16'b0000000000000100: out_v[251] = 10'b1101101100;
    16'b0000000001000100: out_v[251] = 10'b1001001110;
    16'b0000001011000101: out_v[251] = 10'b1010111001;
    16'b0000000000100101: out_v[251] = 10'b1101010111;
    16'b0000100000100100: out_v[251] = 10'b0110001010;
    16'b0000000001000001: out_v[251] = 10'b1010110100;
    16'b0000000001000101: out_v[251] = 10'b1001111010;
    16'b0000100000000100: out_v[251] = 10'b1110001110;
    16'b0000000001100100: out_v[251] = 10'b0011100111;
    16'b0000000000000001: out_v[251] = 10'b1100100011;
    16'b0000000001100000: out_v[251] = 10'b0110010010;
    16'b0000001011000001: out_v[251] = 10'b0101100111;
    16'b0000000000000101: out_v[251] = 10'b0111011011;
    16'b0000001010000001: out_v[251] = 10'b0101001110;
    16'b0000001010000101: out_v[251] = 10'b0111101111;
    16'b0000100000100000: out_v[251] = 10'b0100011010;
    16'b0000101010000001: out_v[251] = 10'b0110110011;
    16'b0000100000000001: out_v[251] = 10'b0000110111;
    16'b0000100000110100: out_v[251] = 10'b0101111000;
    16'b0000100001100000: out_v[251] = 10'b1100110000;
    16'b0000101011100001: out_v[251] = 10'b0011011011;
    16'b0000101011000001: out_v[251] = 10'b0011001010;
    16'b0000101011000000: out_v[251] = 10'b1011101101;
    16'b0000101001000000: out_v[251] = 10'b1100111101;
    16'b0000100000110000: out_v[251] = 10'b1111001000;
    16'b0000100001000100: out_v[251] = 10'b1111010110;
    16'b0000100011000001: out_v[251] = 10'b0101110010;
    16'b0000100001100100: out_v[251] = 10'b1011100111;
    16'b0000000000111000: out_v[251] = 10'b1001000111;
    16'b0000100000011000: out_v[251] = 10'b0011010101;
    16'b0000000000101000: out_v[251] = 10'b1111000011;
    16'b0000100000010100: out_v[251] = 10'b1101011010;
    16'b0100000000000000: out_v[251] = 10'b0101011100;
    16'b0100000000010000: out_v[251] = 10'b1000110011;
    default: out_v[251] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001000000000010: out_v[252] = 10'b0111101001;
    16'b0001000010000000: out_v[252] = 10'b0010111011;
    16'b0001000011010000: out_v[252] = 10'b0110100101;
    16'b0000000010000000: out_v[252] = 10'b0010000101;
    16'b0001000000000000: out_v[252] = 10'b0010110011;
    16'b0001000010010000: out_v[252] = 10'b0101111111;
    16'b0000000000000000: out_v[252] = 10'b1111010111;
    16'b0010000010000000: out_v[252] = 10'b1011111000;
    16'b0011000000000000: out_v[252] = 10'b1000011000;
    16'b0000000010010010: out_v[252] = 10'b1001110111;
    16'b0000000010000010: out_v[252] = 10'b1100110100;
    16'b0001000010000010: out_v[252] = 10'b0011010111;
    16'b0011000010000000: out_v[252] = 10'b1010011101;
    16'b0000000010010100: out_v[252] = 10'b0011111111;
    16'b0000000000000010: out_v[252] = 10'b0111101000;
    16'b0000000010010000: out_v[252] = 10'b0100100111;
    16'b0000000010000100: out_v[252] = 10'b1000110100;
    16'b0000000011010000: out_v[252] = 10'b0111000111;
    16'b0001000011010100: out_v[252] = 10'b1100010111;
    16'b0001000010010100: out_v[252] = 10'b1100101011;
    16'b1001000011010100: out_v[252] = 10'b1010000001;
    16'b0001000010000100: out_v[252] = 10'b0111011000;
    16'b0001000010010010: out_v[252] = 10'b0111110111;
    16'b0010000000000010: out_v[252] = 10'b0110100100;
    16'b0010000000000000: out_v[252] = 10'b1101000110;
    16'b0011000000000010: out_v[252] = 10'b0110101010;
    16'b0010000000000100: out_v[252] = 10'b0101001001;
    16'b1010000000000100: out_v[252] = 10'b0111100101;
    16'b0011000010000100: out_v[252] = 10'b0001100111;
    16'b0011000000000100: out_v[252] = 10'b0101000011;
    16'b0010000010000100: out_v[252] = 10'b1010001110;
    16'b0001000000000100: out_v[252] = 10'b1011010100;
    16'b1011000000000100: out_v[252] = 10'b0101010000;
    16'b0000000000000100: out_v[252] = 10'b1000001100;
    16'b1001000000000000: out_v[252] = 10'b0011001110;
    16'b1000000000000000: out_v[252] = 10'b1001001110;
    16'b1010000000000000: out_v[252] = 10'b0011001111;
    16'b0010000000010000: out_v[252] = 10'b0011110011;
    16'b1011000000000000: out_v[252] = 10'b1000011111;
    16'b1000000000000100: out_v[252] = 10'b0100111110;
    16'b1001000000000100: out_v[252] = 10'b1100000110;
    16'b0010000000000110: out_v[252] = 10'b0110101000;
    16'b0010000010000110: out_v[252] = 10'b0000100100;
    16'b0000000000000110: out_v[252] = 10'b0110110100;
    16'b1010000010000110: out_v[252] = 10'b0011111101;
    16'b0011000000000110: out_v[252] = 10'b1101110110;
    16'b0011000010000110: out_v[252] = 10'b1000001110;
    16'b0011000010000010: out_v[252] = 10'b0101011011;
    16'b1011000010000110: out_v[252] = 10'b1000011011;
    16'b0010000010000010: out_v[252] = 10'b0110110001;
    16'b1011000010000100: out_v[252] = 10'b0010011111;
    16'b1010000010000100: out_v[252] = 10'b0000110010;
    16'b0011000001010000: out_v[252] = 10'b1011111100;
    16'b0011000000010000: out_v[252] = 10'b1010001000;
    16'b0000000000010000: out_v[252] = 10'b1101010111;
    16'b0001000000010000: out_v[252] = 10'b0110100101;
    16'b0001000000000001: out_v[252] = 10'b1100101111;
    16'b0010000010010000: out_v[252] = 10'b0011101110;
    16'b0000010000000000: out_v[252] = 10'b1110100110;
    16'b0010000010100000: out_v[252] = 10'b0000000011;
    16'b0010000010010100: out_v[252] = 10'b0101110101;
    16'b0010000000100000: out_v[252] = 10'b1101101011;
    16'b0000000010100000: out_v[252] = 10'b0011100000;
    16'b0000000000100000: out_v[252] = 10'b1111101100;
    16'b0010010000000000: out_v[252] = 10'b0111100001;
    16'b0010000000010100: out_v[252] = 10'b0011011011;
    16'b0001000001010000: out_v[252] = 10'b0100011101;
    16'b0001001000010010: out_v[252] = 10'b1100111011;
    16'b0010000001010000: out_v[252] = 10'b1101100111;
    16'b0001001000000010: out_v[252] = 10'b1111100100;
    16'b0011001000000010: out_v[252] = 10'b1101001110;
    16'b0011000001010010: out_v[252] = 10'b1001011101;
    16'b0011001001010010: out_v[252] = 10'b0100011100;
    16'b0000001000000010: out_v[252] = 10'b1110000101;
    16'b0001000000010010: out_v[252] = 10'b0011110110;
    16'b0001001001010010: out_v[252] = 10'b0111010000;
    16'b0001001000000000: out_v[252] = 10'b1001010111;
    16'b0000000001010000: out_v[252] = 10'b1001011000;
    16'b0011001000000000: out_v[252] = 10'b1110001101;
    16'b0001000001010010: out_v[252] = 10'b0011111011;
    16'b0011001000010010: out_v[252] = 10'b1101111111;
    16'b0011000000010010: out_v[252] = 10'b1101100110;
    16'b0010001000000010: out_v[252] = 10'b1110000001;
    16'b0010000000010010: out_v[252] = 10'b1001011011;
    default: out_v[252] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010000000100001: out_v[253] = 10'b1000100010;
    16'b1011100100000001: out_v[253] = 10'b0011011001;
    16'b1010100000000000: out_v[253] = 10'b0101000011;
    16'b1010000000100001: out_v[253] = 10'b1000110101;
    16'b1011100000100001: out_v[253] = 10'b0000010101;
    16'b1010100000100000: out_v[253] = 10'b1111100001;
    16'b1000100000000000: out_v[253] = 10'b0010000101;
    16'b1010000000000001: out_v[253] = 10'b1001010110;
    16'b1011100000000000: out_v[253] = 10'b0110011010;
    16'b1000000000000000: out_v[253] = 10'b0000011111;
    16'b1011100000000001: out_v[253] = 10'b0001110011;
    16'b1010100000100001: out_v[253] = 10'b1001101111;
    16'b1010100000000001: out_v[253] = 10'b0111100110;
    16'b1010100010100001: out_v[253] = 10'b1001101011;
    16'b0010000000000001: out_v[253] = 10'b0011110100;
    16'b0010100000100000: out_v[253] = 10'b0001011111;
    16'b1000000000100000: out_v[253] = 10'b0011001010;
    16'b1000100000100000: out_v[253] = 10'b0001111011;
    16'b0000000010000000: out_v[253] = 10'b1110110011;
    16'b1000000010000000: out_v[253] = 10'b1110110000;
    16'b1010100010100000: out_v[253] = 10'b1011100011;
    16'b0000100010000000: out_v[253] = 10'b1101100101;
    16'b1001100000000000: out_v[253] = 10'b1001001011;
    16'b1000000010100000: out_v[253] = 10'b1110100011;
    16'b1010000000000000: out_v[253] = 10'b0001110100;
    16'b1010000000100000: out_v[253] = 10'b1100100001;
    16'b0000100010100000: out_v[253] = 10'b1111010101;
    16'b0000000000000000: out_v[253] = 10'b1000010010;
    16'b0000000000100000: out_v[253] = 10'b0000000110;
    16'b1000100010100000: out_v[253] = 10'b0011010111;
    16'b0000100000000000: out_v[253] = 10'b1101100111;
    16'b1000100010000000: out_v[253] = 10'b1101110010;
    16'b0010000000000000: out_v[253] = 10'b1101001010;
    16'b0000000100100000: out_v[253] = 10'b1010101011;
    16'b0001000000100000: out_v[253] = 10'b0001110000;
    16'b0010000000100000: out_v[253] = 10'b0111010101;
    16'b0010000010100000: out_v[253] = 10'b0101100110;
    16'b1000000000100001: out_v[253] = 10'b0001011100;
    16'b0010000010000001: out_v[253] = 10'b0011101110;
    16'b0010100000100001: out_v[253] = 10'b1011000110;
    16'b0000000010100000: out_v[253] = 10'b0001110101;
    16'b0010000010100001: out_v[253] = 10'b1000100110;
    16'b0000000000100001: out_v[253] = 10'b1100001010;
    16'b0000000000000001: out_v[253] = 10'b0010111001;
    16'b0010000100000000: out_v[253] = 10'b0110011011;
    16'b0000000010000001: out_v[253] = 10'b0111100011;
    16'b0010000100000001: out_v[253] = 10'b1010100110;
    16'b1000000010000001: out_v[253] = 10'b1101100101;
    16'b0010000010000000: out_v[253] = 10'b0111011011;
    16'b1010000100000001: out_v[253] = 10'b0001111001;
    16'b0000000100000001: out_v[253] = 10'b1001001110;
    16'b1000000000000001: out_v[253] = 10'b0101011000;
    16'b0000000100000000: out_v[253] = 10'b1101001100;
    16'b0010000110000001: out_v[253] = 10'b1101011010;
    16'b1010000010000001: out_v[253] = 10'b1001111110;
    16'b1010000010000000: out_v[253] = 10'b0111110010;
    16'b1001000000000001: out_v[253] = 10'b1111100100;
    16'b1001000000000000: out_v[253] = 10'b1000111111;
    16'b1001000000100000: out_v[253] = 10'b1001010000;
    16'b1001000000100001: out_v[253] = 10'b0000011001;
    16'b1011000000000001: out_v[253] = 10'b1011100110;
    16'b1010000010000011: out_v[253] = 10'b0010010111;
    16'b1010000010100001: out_v[253] = 10'b1001001011;
    16'b1011000000100001: out_v[253] = 10'b1101011000;
    16'b0001000000000000: out_v[253] = 10'b1100010100;
    16'b0011000000000001: out_v[253] = 10'b0111100010;
    16'b0011000000000000: out_v[253] = 10'b1100100010;
    16'b1011000000000000: out_v[253] = 10'b0110100100;
    16'b0011000000100001: out_v[253] = 10'b0100001010;
    16'b1011000000100000: out_v[253] = 10'b0100110010;
    16'b0011000000100000: out_v[253] = 10'b1100000111;
    16'b0000100000100000: out_v[253] = 10'b1100010010;
    16'b1011000100000001: out_v[253] = 10'b0111111010;
    16'b0011000100000001: out_v[253] = 10'b0010110111;
    16'b1010000010100000: out_v[253] = 10'b0111001001;
    16'b0010001000000011: out_v[253] = 10'b1101110100;
    16'b0010000010000011: out_v[253] = 10'b0011100010;
    16'b0010001010000001: out_v[253] = 10'b0000111110;
    16'b0010001010000011: out_v[253] = 10'b0111100101;
    16'b1010001000000001: out_v[253] = 10'b0000010011;
    16'b0000001000000000: out_v[253] = 10'b1100100001;
    16'b0010001010000000: out_v[253] = 10'b1101111111;
    16'b0010001000000001: out_v[253] = 10'b1001001111;
    16'b0000001010000000: out_v[253] = 10'b0111011001;
    16'b0001000100100000: out_v[253] = 10'b1101000011;
    16'b1010001010000001: out_v[253] = 10'b0110100110;
    16'b0010001000000000: out_v[253] = 10'b0011001111;
    16'b0010000000000011: out_v[253] = 10'b1111101011;
    16'b0010000100100001: out_v[253] = 10'b1001111011;
    16'b1010001000000000: out_v[253] = 10'b0011000011;
    16'b0001000100000000: out_v[253] = 10'b0111011111;
    16'b0001100000100000: out_v[253] = 10'b1011000100;
    16'b0000000010100001: out_v[253] = 10'b1100010011;
    16'b1000000010100001: out_v[253] = 10'b0101100110;
    16'b0001100100100000: out_v[253] = 10'b0011101111;
    16'b1000001000000000: out_v[253] = 10'b1100101111;
    default: out_v[253] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000010100001010: out_v[254] = 10'b0100110011;
    16'b1010110000001010: out_v[254] = 10'b1101100100;
    16'b1100010100000010: out_v[254] = 10'b0111011011;
    16'b0100010100000010: out_v[254] = 10'b1100011011;
    16'b0010010000001010: out_v[254] = 10'b1001000101;
    16'b1000010000001000: out_v[254] = 10'b0111001011;
    16'b1010010000000010: out_v[254] = 10'b0000110101;
    16'b0110000100001010: out_v[254] = 10'b0110110011;
    16'b1000110000001010: out_v[254] = 10'b0010110000;
    16'b1010010000001010: out_v[254] = 10'b1100111110;
    16'b0110110000001010: out_v[254] = 10'b1011110010;
    16'b1010010100001010: out_v[254] = 10'b1111010110;
    16'b1110010110001010: out_v[254] = 10'b1110101011;
    16'b0110010100001010: out_v[254] = 10'b0011111010;
    16'b1110010100001010: out_v[254] = 10'b1000010010;
    16'b1100010100001010: out_v[254] = 10'b0011111110;
    16'b1100010100001000: out_v[254] = 10'b1101101100;
    16'b1100010110001010: out_v[254] = 10'b1011111110;
    16'b1000010110001000: out_v[254] = 10'b1101100111;
    16'b1000010110001010: out_v[254] = 10'b1010111111;
    16'b1000010100001000: out_v[254] = 10'b0100010101;
    16'b1000010100001010: out_v[254] = 10'b1011001011;
    16'b1100010110000000: out_v[254] = 10'b0111001011;
    16'b0110010000001010: out_v[254] = 10'b0111110011;
    16'b0010110000001000: out_v[254] = 10'b0000111011;
    16'b0110010100000010: out_v[254] = 10'b1011001111;
    16'b1010011000101010: out_v[254] = 10'b0111111010;
    16'b1010000000001010: out_v[254] = 10'b0001011011;
    16'b1100010110000010: out_v[254] = 10'b1100110101;
    16'b1010111000101010: out_v[254] = 10'b1111110011;
    16'b1000010000000000: out_v[254] = 10'b1111001001;
    16'b0010111000001010: out_v[254] = 10'b0100010111;
    16'b1000010100000000: out_v[254] = 10'b1010110010;
    16'b0010110000001010: out_v[254] = 10'b1000111100;
    16'b1010110000000010: out_v[254] = 10'b0010011111;
    16'b0010010100001010: out_v[254] = 10'b0011100010;
    16'b1000010000001010: out_v[254] = 10'b1011000000;
    16'b0110010000000010: out_v[254] = 10'b0100010011;
    16'b1100010100000000: out_v[254] = 10'b0010101011;
    16'b1010010000101010: out_v[254] = 10'b0010101011;
    16'b1110110000001010: out_v[254] = 10'b1011111011;
    16'b1100010110001000: out_v[254] = 10'b1000110001;
    16'b1000110100001010: out_v[254] = 10'b1111000001;
    16'b1110010000001010: out_v[254] = 10'b1111110110;
    16'b1000000000001010: out_v[254] = 10'b0010111011;
    16'b1000010100000010: out_v[254] = 10'b1101001111;
    16'b1100010000001010: out_v[254] = 10'b1100111110;
    16'b1010110000101010: out_v[254] = 10'b1111011011;
    16'b1110110100001010: out_v[254] = 10'b1001111111;
    16'b1110010100000010: out_v[254] = 10'b0110000011;
    16'b1010110100001010: out_v[254] = 10'b1000101111;
    16'b0000100000001000: out_v[254] = 10'b1001000011;
    16'b0000010000000000: out_v[254] = 10'b0111100111;
    16'b0000100000000000: out_v[254] = 10'b0111010000;
    16'b0000100100000000: out_v[254] = 10'b1110001010;
    16'b0100100000000000: out_v[254] = 10'b1110011010;
    16'b0100100000001000: out_v[254] = 10'b1011000110;
    16'b0000000000001000: out_v[254] = 10'b1011100111;
    16'b0100100100000000: out_v[254] = 10'b1100100110;
    16'b0010100100000000: out_v[254] = 10'b0101011011;
    16'b0000000000000000: out_v[254] = 10'b0100001110;
    16'b0000100110000000: out_v[254] = 10'b0110000000;
    16'b0010100110000000: out_v[254] = 10'b1110001011;
    16'b0000011000000000: out_v[254] = 10'b0111100010;
    16'b0000110000000000: out_v[254] = 10'b0111110000;
    16'b0100000000001000: out_v[254] = 10'b1100110011;
    16'b0000111000000000: out_v[254] = 10'b0010000111;
    16'b0000110000001000: out_v[254] = 10'b1101010000;
    16'b0100000000000000: out_v[254] = 10'b1101010100;
    16'b0000000110001000: out_v[254] = 10'b1011111001;
    16'b0100100110001000: out_v[254] = 10'b1101001100;
    16'b0010000110001000: out_v[254] = 10'b1001011010;
    16'b0100000110001000: out_v[254] = 10'b1011011100;
    16'b0000000100001000: out_v[254] = 10'b0011101101;
    16'b0010000000000000: out_v[254] = 10'b1001110001;
    16'b0110010000000000: out_v[254] = 10'b0010110110;
    16'b0100000110000000: out_v[254] = 10'b1001100011;
    16'b0110000110001000: out_v[254] = 10'b1001100100;
    16'b0110000010001000: out_v[254] = 10'b0101010111;
    16'b0110000110000000: out_v[254] = 10'b1010111010;
    16'b0110010010000000: out_v[254] = 10'b1110000111;
    16'b0010000000001000: out_v[254] = 10'b0010110000;
    16'b0100000010001000: out_v[254] = 10'b1111100000;
    16'b0110011100000000: out_v[254] = 10'b1101110110;
    16'b0110010100000000: out_v[254] = 10'b1110101100;
    16'b0110010110100000: out_v[254] = 10'b1101001011;
    16'b0100000100000000: out_v[254] = 10'b1001010111;
    16'b0100000010000000: out_v[254] = 10'b1011111100;
    16'b0110000010000000: out_v[254] = 10'b0110000011;
    16'b0110000100000000: out_v[254] = 10'b1101100111;
    16'b0010000100001000: out_v[254] = 10'b0111100101;
    16'b0110010110001000: out_v[254] = 10'b0111011011;
    16'b0100010100000000: out_v[254] = 10'b1011001111;
    16'b0100010010000000: out_v[254] = 10'b1010110101;
    16'b0010010000001000: out_v[254] = 10'b1011011010;
    16'b0110010100100000: out_v[254] = 10'b1010101110;
    16'b0010000110000000: out_v[254] = 10'b1001000100;
    16'b0010010100001000: out_v[254] = 10'b0111101011;
    16'b0100000100001000: out_v[254] = 10'b1001010011;
    16'b0110000100001000: out_v[254] = 10'b0010011111;
    16'b0110010110000000: out_v[254] = 10'b1100110001;
    16'b0010100000000000: out_v[254] = 10'b0011010100;
    16'b0100100010001000: out_v[254] = 10'b0111011100;
    16'b0110010100001000: out_v[254] = 10'b1011110110;
    16'b0010000010001000: out_v[254] = 10'b1000100111;
    16'b0010010000101000: out_v[254] = 10'b1001100110;
    16'b0000010100001000: out_v[254] = 10'b0000101111;
    16'b0100010110000000: out_v[254] = 10'b0011111111;
    16'b0010000100000000: out_v[254] = 10'b1111000111;
    16'b0110010000100000: out_v[254] = 10'b0111110011;
    16'b0110100110001000: out_v[254] = 10'b1110100001;
    16'b0010101100001000: out_v[254] = 10'b1110110111;
    16'b0110100100000000: out_v[254] = 10'b1100100001;
    16'b0010100100000010: out_v[254] = 10'b1010010101;
    16'b0000100100001000: out_v[254] = 10'b1100111100;
    16'b0010100100001000: out_v[254] = 10'b0001010101;
    16'b0010111100101010: out_v[254] = 10'b1011111110;
    16'b1000100100001010: out_v[254] = 10'b0000101010;
    16'b0000100100001010: out_v[254] = 10'b0111110010;
    16'b0110100010000000: out_v[254] = 10'b0110111001;
    16'b0110100100001000: out_v[254] = 10'b0111011010;
    16'b0110100000001000: out_v[254] = 10'b1000001101;
    16'b0010110100001010: out_v[254] = 10'b1001101110;
    16'b0010100100001010: out_v[254] = 10'b1000101100;
    16'b0010110100001000: out_v[254] = 10'b0101010011;
    16'b0000100100000010: out_v[254] = 10'b0001111000;
    16'b0010100000001000: out_v[254] = 10'b1001110001;
    16'b0010111100101000: out_v[254] = 10'b0100110011;
    16'b0100100110001010: out_v[254] = 10'b1000011110;
    16'b0010111100001010: out_v[254] = 10'b0011001111;
    16'b0010100110001010: out_v[254] = 10'b0011101111;
    16'b0010100110001000: out_v[254] = 10'b1011111001;
    16'b0000110100001000: out_v[254] = 10'b0111000000;
    16'b0000100110001010: out_v[254] = 10'b0111110111;
    16'b0110100110001010: out_v[254] = 10'b1111001110;
    16'b0100100010001010: out_v[254] = 10'b1000001100;
    16'b0010011100001000: out_v[254] = 10'b0011111100;
    16'b0010111100001000: out_v[254] = 10'b0100010100;
    16'b0110100110000000: out_v[254] = 10'b0010110011;
    16'b0110100010001000: out_v[254] = 10'b0010111011;
    16'b0010000000000010: out_v[254] = 10'b0100110001;
    16'b0010000000001010: out_v[254] = 10'b0010110100;
    16'b0010010100000010: out_v[254] = 10'b0001110000;
    16'b1000000000000010: out_v[254] = 10'b0001011011;
    16'b0010000100000010: out_v[254] = 10'b1000011110;
    16'b0010110000000010: out_v[254] = 10'b0010110010;
    16'b0010010000000010: out_v[254] = 10'b0100110010;
    16'b0010010000000000: out_v[254] = 10'b1101010100;
    16'b0000010100000010: out_v[254] = 10'b1101000011;
    16'b0000000000001010: out_v[254] = 10'b1011000011;
    16'b0000000000000010: out_v[254] = 10'b0101010001;
    16'b0000110000000010: out_v[254] = 10'b0010100101;
    16'b0010000100001010: out_v[254] = 10'b1010000111;
    16'b0010110100000010: out_v[254] = 10'b0101110110;
    16'b1010000000000010: out_v[254] = 10'b1110101011;
    16'b0010100000000010: out_v[254] = 10'b1011000101;
    16'b0000010000000010: out_v[254] = 10'b0101101000;
    16'b0110000000001010: out_v[254] = 10'b0110010011;
    16'b1010010000000000: out_v[254] = 10'b0001011110;
    16'b0010100000001010: out_v[254] = 10'b0111111110;
    16'b1010010100000010: out_v[254] = 10'b0100110100;
    16'b0010010110000010: out_v[254] = 10'b0111111011;
    16'b1000010000000010: out_v[254] = 10'b1010111111;
    16'b0010010100000000: out_v[254] = 10'b1011101110;
    16'b1010100000001010: out_v[254] = 10'b1001110010;
    16'b0010110000000000: out_v[254] = 10'b0110100010;
    16'b0000000100001010: out_v[254] = 10'b1110100001;
    16'b0000000100000010: out_v[254] = 10'b1000100111;
    16'b0000100000001010: out_v[254] = 10'b1001110000;
    16'b0000010000001010: out_v[254] = 10'b1000100111;
    16'b0000100000000010: out_v[254] = 10'b1100101110;
    16'b0100100100000010: out_v[254] = 10'b1111010010;
    16'b0100100110000010: out_v[254] = 10'b1010100111;
    16'b0110100100000010: out_v[254] = 10'b0011111100;
    16'b0110100000001010: out_v[254] = 10'b1011000111;
    16'b0110000000000010: out_v[254] = 10'b0111111001;
    16'b1010000010000010: out_v[254] = 10'b1110100111;
    16'b0110100000000010: out_v[254] = 10'b1000100111;
    16'b1010000110000010: out_v[254] = 10'b1001001110;
    16'b1110000110000010: out_v[254] = 10'b1111001000;
    16'b0110100000000000: out_v[254] = 10'b1011000000;
    16'b1100000100000010: out_v[254] = 10'b1011101000;
    16'b1110000100000010: out_v[254] = 10'b0110111010;
    16'b0100000100000010: out_v[254] = 10'b0010001111;
    16'b1000000010000010: out_v[254] = 10'b0011111010;
    16'b1110000000000010: out_v[254] = 10'b1001100100;
    16'b1100000110000010: out_v[254] = 10'b0001100111;
    16'b0110000100000010: out_v[254] = 10'b1111001111;
    16'b1100000000000010: out_v[254] = 10'b0111000011;
    16'b1110100100000010: out_v[254] = 10'b1110110011;
    16'b0110000000000000: out_v[254] = 10'b0000011110;
    16'b0010000110000010: out_v[254] = 10'b0110111001;
    16'b0100000000000010: out_v[254] = 10'b1101101011;
    16'b1000000110000010: out_v[254] = 10'b1110010111;
    16'b0000000110000010: out_v[254] = 10'b1010011111;
    16'b1100100100000010: out_v[254] = 10'b1101010010;
    16'b0110000110000010: out_v[254] = 10'b0110100011;
    16'b1110100000001010: out_v[254] = 10'b1110100110;
    16'b0000010000001000: out_v[254] = 10'b0011011111;
    16'b0000000100000000: out_v[254] = 10'b1110011101;
    16'b0110110100000000: out_v[254] = 10'b1100010111;
    16'b0100110000000000: out_v[254] = 10'b0110001000;
    16'b0100110100000000: out_v[254] = 10'b0111001011;
    16'b0000110100001010: out_v[254] = 10'b0010001111;
    16'b0000111000001000: out_v[254] = 10'b1101101000;
    16'b0010110100000000: out_v[254] = 10'b0110010001;
    16'b0000110100000000: out_v[254] = 10'b1101000001;
    16'b0010111000001000: out_v[254] = 10'b0001001111;
    16'b0000010100000000: out_v[254] = 10'b0010000101;
    16'b0000110000001010: out_v[254] = 10'b0000111110;
    default: out_v[254] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000110000000000: out_v[255] = 10'b1101000110;
    16'b0000000000000000: out_v[255] = 10'b0110100010;
    16'b0000001000000000: out_v[255] = 10'b0000110001;
    16'b0000001001000000: out_v[255] = 10'b1110000101;
    16'b0000010000000000: out_v[255] = 10'b0111100101;
    16'b0000011001010000: out_v[255] = 10'b0001000001;
    16'b0000011000000000: out_v[255] = 10'b1001010001;
    16'b0000001001010000: out_v[255] = 10'b0101101001;
    16'b0000011001000000: out_v[255] = 10'b1010110111;
    16'b0000000001010000: out_v[255] = 10'b1111001010;
    16'b0000000001000000: out_v[255] = 10'b1101101110;
    16'b0000101001010000: out_v[255] = 10'b0010101010;
    16'b0000101001000000: out_v[255] = 10'b0100000011;
    16'b0000010001010000: out_v[255] = 10'b0010011100;
    16'b0000100000000000: out_v[255] = 10'b1111100001;
    16'b0000101000000000: out_v[255] = 10'b0010110000;
    16'b0000010001000000: out_v[255] = 10'b1000001101;
    16'b0000010000000100: out_v[255] = 10'b1011100100;
    16'b0000010100000000: out_v[255] = 10'b0000100000;
    16'b0000010000000010: out_v[255] = 10'b1011001101;
    16'b0000010000010000: out_v[255] = 10'b1000001111;
    16'b0000000000010000: out_v[255] = 10'b0111001100;
    16'b0000010100000100: out_v[255] = 10'b0101010100;
    16'b0000000100000000: out_v[255] = 10'b0001001111;
    16'b0000000100000100: out_v[255] = 10'b0011011110;
    16'b0000000000000100: out_v[255] = 10'b0101111010;
    16'b0000100001000000: out_v[255] = 10'b1011111010;
    16'b0010000000000100: out_v[255] = 10'b0100001011;
    16'b1000001000000000: out_v[255] = 10'b1100010100;
    16'b0000000000000001: out_v[255] = 10'b0111110000;
    16'b0000010000000001: out_v[255] = 10'b1011100010;
    16'b0000011000000001: out_v[255] = 10'b0111010010;
    16'b1000100000000000: out_v[255] = 10'b0110111000;
    16'b1000000000000000: out_v[255] = 10'b0110001010;
    16'b1100100000000000: out_v[255] = 10'b0011101010;
    16'b0100100000000000: out_v[255] = 10'b1100010111;
    16'b0000111000000000: out_v[255] = 10'b1100000000;
    default: out_v[255] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000001000101100: out_v[256] = 10'b0010100110;
    16'b0000001000101001: out_v[256] = 10'b1101110001;
    16'b0000000000101000: out_v[256] = 10'b1011100101;
    16'b0101101000101000: out_v[256] = 10'b0010010011;
    16'b0100001000101100: out_v[256] = 10'b1000100001;
    16'b0001101000000000: out_v[256] = 10'b0101100110;
    16'b0100000000101000: out_v[256] = 10'b0111100100;
    16'b0000001000001100: out_v[256] = 10'b0100011111;
    16'b0101001000100000: out_v[256] = 10'b1011001101;
    16'b0001001000101100: out_v[256] = 10'b1111011111;
    16'b0001001000100000: out_v[256] = 10'b0101001010;
    16'b0000001000101000: out_v[256] = 10'b1010110110;
    16'b0100001000101000: out_v[256] = 10'b0110000110;
    16'b0001001000101000: out_v[256] = 10'b1000011000;
    16'b0001001000101001: out_v[256] = 10'b1001011101;
    16'b0100000000101100: out_v[256] = 10'b1001101100;
    16'b0101101000101100: out_v[256] = 10'b0010011010;
    16'b0000000100101000: out_v[256] = 10'b0011011000;
    16'b0000001000001000: out_v[256] = 10'b1101011111;
    16'b0001001000100100: out_v[256] = 10'b1111000100;
    16'b0001101000100001: out_v[256] = 10'b0011001011;
    16'b0001100000000000: out_v[256] = 10'b1010110011;
    16'b0001101000101001: out_v[256] = 10'b0101111100;
    16'b0001101000000001: out_v[256] = 10'b1101110010;
    16'b0000000000100000: out_v[256] = 10'b1110110001;
    16'b0000001000100000: out_v[256] = 10'b1101010110;
    16'b0001101000100000: out_v[256] = 10'b1011010110;
    16'b0101101000100100: out_v[256] = 10'b1100100001;
    16'b0101101000100001: out_v[256] = 10'b1011110011;
    16'b0001000000100000: out_v[256] = 10'b0110010110;
    16'b0000000000001100: out_v[256] = 10'b0100011001;
    16'b0101001000101000: out_v[256] = 10'b1011010010;
    16'b0101001000101100: out_v[256] = 10'b1110100000;
    16'b0101101000101001: out_v[256] = 10'b0111001011;
    16'b0101101000100000: out_v[256] = 10'b0010110110;
    16'b0100001000101001: out_v[256] = 10'b0010100111;
    16'b0101101000000000: out_v[256] = 10'b1010000111;
    16'b0100001000000100: out_v[256] = 10'b1001010001;
    16'b0001001000100001: out_v[256] = 10'b1101000110;
    16'b0101101000000001: out_v[256] = 10'b0000100001;
    16'b0000001000000100: out_v[256] = 10'b0100110011;
    16'b0101101000101101: out_v[256] = 10'b1000101011;
    16'b0000000000101100: out_v[256] = 10'b1100000110;
    16'b0101001000101001: out_v[256] = 10'b1111011100;
    16'b0000000000101001: out_v[256] = 10'b0001100010;
    16'b0000000000000100: out_v[256] = 10'b1111001100;
    16'b0000001000000000: out_v[256] = 10'b1000111010;
    16'b0001000000101000: out_v[256] = 10'b0001011110;
    16'b0101000000001100: out_v[256] = 10'b0011100110;
    16'b0100000000000000: out_v[256] = 10'b0101000111;
    16'b0000000000000000: out_v[256] = 10'b1010111100;
    16'b0001000000000100: out_v[256] = 10'b1100000010;
    16'b0100000000001100: out_v[256] = 10'b0011111011;
    16'b0100000000000100: out_v[256] = 10'b1010000101;
    16'b0101000000101100: out_v[256] = 10'b0011011010;
    16'b0100000000001000: out_v[256] = 10'b1101010101;
    16'b0101000000000100: out_v[256] = 10'b1101001100;
    16'b0001100000101101: out_v[256] = 10'b1010110111;
    16'b0001100000101100: out_v[256] = 10'b0010110110;
    16'b0101100000101100: out_v[256] = 10'b0000011011;
    16'b0110000000000000: out_v[256] = 10'b0011000010;
    16'b0001000000001100: out_v[256] = 10'b1111100000;
    16'b0001000000101100: out_v[256] = 10'b0010010011;
    16'b0100000100000100: out_v[256] = 10'b1000101100;
    16'b0100000100101100: out_v[256] = 10'b0111110110;
    16'b0110000000001100: out_v[256] = 10'b1000111111;
    16'b0000000100001100: out_v[256] = 10'b1010110111;
    16'b0101100000100101: out_v[256] = 10'b1001010100;
    16'b0100000000101101: out_v[256] = 10'b1010110001;
    16'b0000000100000100: out_v[256] = 10'b0100100110;
    16'b0110000000101100: out_v[256] = 10'b1010101100;
    16'b0101000000101101: out_v[256] = 10'b0001100011;
    16'b0000000100101100: out_v[256] = 10'b1110000100;
    16'b0100000100001100: out_v[256] = 10'b1101011010;
    16'b0110000000000100: out_v[256] = 10'b1011100101;
    16'b0100000100000000: out_v[256] = 10'b1100010101;
    16'b0111000000101100: out_v[256] = 10'b0110010101;
    16'b0100000000101001: out_v[256] = 10'b1011111100;
    16'b0101100000101101: out_v[256] = 10'b1100000101;
    16'b0111100000101101: out_v[256] = 10'b0111111011;
    16'b1100000000000100: out_v[256] = 10'b0101101100;
    16'b0100000100101000: out_v[256] = 10'b0101111111;
    16'b1100000100000100: out_v[256] = 10'b0111011010;
    16'b1000000000000100: out_v[256] = 10'b1101000110;
    16'b0111000000101101: out_v[256] = 10'b1011000111;
    16'b0110000000101101: out_v[256] = 10'b1111100011;
    16'b0000000000000001: out_v[256] = 10'b0101111101;
    16'b0000001100000000: out_v[256] = 10'b0000111010;
    16'b0101100000101001: out_v[256] = 10'b0001011111;
    16'b0000000000001000: out_v[256] = 10'b1011011001;
    16'b0000001100000001: out_v[256] = 10'b1011110111;
    16'b0101000000101001: out_v[256] = 10'b1011100111;
    16'b0001100000101001: out_v[256] = 10'b1111011001;
    16'b0101000000101000: out_v[256] = 10'b0100011011;
    16'b0000001000001001: out_v[256] = 10'b0111001111;
    16'b0001000000101001: out_v[256] = 10'b1000011011;
    16'b0000000100000001: out_v[256] = 10'b0110001010;
    16'b0100001000000000: out_v[256] = 10'b0111011100;
    16'b0000000100000000: out_v[256] = 10'b1000011011;
    16'b0000000100001000: out_v[256] = 10'b1010001111;
    16'b0000001000000001: out_v[256] = 10'b1011100101;
    16'b0000000000001001: out_v[256] = 10'b0100110111;
    16'b0100001000001100: out_v[256] = 10'b1100010001;
    16'b0100001000100000: out_v[256] = 10'b0110110111;
    16'b0001101000101100: out_v[256] = 10'b0101100101;
    16'b0101001000001100: out_v[256] = 10'b1000110011;
    16'b0100101000100000: out_v[256] = 10'b1101101111;
    16'b0100001000100100: out_v[256] = 10'b0000110010;
    16'b0001101000101000: out_v[256] = 10'b0001101100;
    16'b0100001000001000: out_v[256] = 10'b0111001111;
    16'b0001101000100100: out_v[256] = 10'b0111001011;
    16'b0001001000000000: out_v[256] = 10'b0100100010;
    16'b0001000000000000: out_v[256] = 10'b0011110101;
    16'b0101100000000000: out_v[256] = 10'b0010100001;
    16'b0101100000000100: out_v[256] = 10'b1111101010;
    16'b0101101000000100: out_v[256] = 10'b1100001001;
    16'b0001100000000001: out_v[256] = 10'b1011100001;
    16'b0001101000000100: out_v[256] = 10'b0001000101;
    16'b0001001000000100: out_v[256] = 10'b1001001110;
    16'b0101100000101000: out_v[256] = 10'b1100100001;
    16'b0001100000000100: out_v[256] = 10'b1011110111;
    16'b0110001000000100: out_v[256] = 10'b0111101000;
    16'b0100001100000100: out_v[256] = 10'b0011001011;
    16'b0110001000000000: out_v[256] = 10'b0011101000;
    16'b0100001100101100: out_v[256] = 10'b1011001110;
    16'b0100001001000100: out_v[256] = 10'b0001100011;
    16'b0010000000000100: out_v[256] = 10'b1101011000;
    16'b0010001000000100: out_v[256] = 10'b1011001010;
    16'b0101001000000100: out_v[256] = 10'b1111101001;
    16'b0000010000101000: out_v[256] = 10'b0101011011;
    16'b0000010000010000: out_v[256] = 10'b1010100010;
    16'b0000000000111000: out_v[256] = 10'b1001100101;
    16'b0100000000111000: out_v[256] = 10'b0110110110;
    16'b0000000000010000: out_v[256] = 10'b1110000011;
    16'b0000010000111000: out_v[256] = 10'b1101111101;
    16'b0100000000100000: out_v[256] = 10'b1101000111;
    16'b0100010000111000: out_v[256] = 10'b0101010001;
    16'b0000001000100100: out_v[256] = 10'b1101000111;
    16'b0101000000100100: out_v[256] = 10'b1110101111;
    16'b0100000000100100: out_v[256] = 10'b0011111000;
    16'b0001000000100100: out_v[256] = 10'b1101011001;
    16'b0101100000100100: out_v[256] = 10'b0100011101;
    16'b0001100000100100: out_v[256] = 10'b1010011101;
    16'b0000000000100100: out_v[256] = 10'b1100000111;
    16'b0101001000100100: out_v[256] = 10'b1100011111;
    default: out_v[256] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000000000000: out_v[257] = 10'b0011010011;
    16'b0000101000001010: out_v[257] = 10'b1100000010;
    16'b0000101000100010: out_v[257] = 10'b0001001001;
    16'b0000101000000010: out_v[257] = 10'b0001001100;
    16'b0000100000000010: out_v[257] = 10'b0000101011;
    16'b0000100000100010: out_v[257] = 10'b1101000111;
    16'b0000100000000000: out_v[257] = 10'b1111010011;
    16'b0000000000100000: out_v[257] = 10'b0111010001;
    16'b0000001000000010: out_v[257] = 10'b0100001101;
    16'b0000001000100010: out_v[257] = 10'b1111000111;
    16'b0000100000100000: out_v[257] = 10'b0011010111;
    16'b0000001000000000: out_v[257] = 10'b0100110000;
    16'b0001100000000010: out_v[257] = 10'b1011011100;
    16'b0000101000000000: out_v[257] = 10'b0100010110;
    16'b0001100000100010: out_v[257] = 10'b1011010011;
    16'b0000000000000010: out_v[257] = 10'b0000000101;
    16'b0000001000001000: out_v[257] = 10'b1011011000;
    16'b0001000000000000: out_v[257] = 10'b1100110110;
    16'b0001101000000010: out_v[257] = 10'b1000110111;
    16'b0001001000000000: out_v[257] = 10'b0000101111;
    16'b0001000000000010: out_v[257] = 10'b1011010110;
    16'b0000000100000000: out_v[257] = 10'b0010010110;
    16'b0001100000000000: out_v[257] = 10'b0111001011;
    16'b0000001010001000: out_v[257] = 10'b0010111100;
    16'b0100001000001000: out_v[257] = 10'b0011001010;
    16'b0100001000000000: out_v[257] = 10'b1011111000;
    16'b0000000010000000: out_v[257] = 10'b0011011011;
    16'b0000001000001010: out_v[257] = 10'b0000101011;
    16'b0000001010000000: out_v[257] = 10'b0000101011;
    16'b0000000000000001: out_v[257] = 10'b1011000000;
    16'b0000000010000001: out_v[257] = 10'b0001110001;
    16'b0000000011000000: out_v[257] = 10'b1001001100;
    16'b0000000000000100: out_v[257] = 10'b0010000001;
    16'b0000001011001000: out_v[257] = 10'b1111000011;
    16'b0000001011000000: out_v[257] = 10'b1100001111;
    default: out_v[257] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010000001100001: out_v[258] = 10'b1000010010;
    16'b0010010011100011: out_v[258] = 10'b1000110110;
    16'b0010000001100010: out_v[258] = 10'b1100101011;
    16'b0010000001100000: out_v[258] = 10'b0110001110;
    16'b0010000001100011: out_v[258] = 10'b1000011011;
    16'b0010000000100010: out_v[258] = 10'b1111001011;
    16'b0010000000100001: out_v[258] = 10'b1001111101;
    16'b0010000001110001: out_v[258] = 10'b0110101110;
    16'b0010000001000001: out_v[258] = 10'b0101011010;
    16'b0000000001100010: out_v[258] = 10'b0010111111;
    16'b0010000001000010: out_v[258] = 10'b0000111110;
    16'b0000000001100011: out_v[258] = 10'b1110000011;
    16'b0010010011100010: out_v[258] = 10'b1100100011;
    16'b0010010001100011: out_v[258] = 10'b0111011010;
    16'b0000000001100001: out_v[258] = 10'b1100110011;
    16'b0011000001100011: out_v[258] = 10'b0100101011;
    16'b0010010010100011: out_v[258] = 10'b0001100100;
    16'b0010010010100010: out_v[258] = 10'b0110110010;
    16'b0010000000100011: out_v[258] = 10'b0011011111;
    16'b0010000011100010: out_v[258] = 10'b0111010011;
    16'b0010000010100010: out_v[258] = 10'b1111001000;
    16'b0010000001000011: out_v[258] = 10'b0101011111;
    16'b0010000000000001: out_v[258] = 10'b1000111111;
    16'b0010000001110011: out_v[258] = 10'b0001011111;
    16'b0010000000100000: out_v[258] = 10'b0011001110;
    16'b0010000001000000: out_v[258] = 10'b0010110111;
    16'b0010010001100010: out_v[258] = 10'b0111100011;
    16'b0010000011100011: out_v[258] = 10'b0010111111;
    16'b0010000000110000: out_v[258] = 10'b0000101100;
    16'b0000000000010000: out_v[258] = 10'b0001011110;
    16'b0000000000010001: out_v[258] = 10'b1111000111;
    16'b0010000000010001: out_v[258] = 10'b1101000110;
    16'b0010000000010000: out_v[258] = 10'b0010100110;
    16'b0000000000110000: out_v[258] = 10'b0001010010;
    16'b0010000000110001: out_v[258] = 10'b1100100000;
    16'b0000000000110001: out_v[258] = 10'b0100110000;
    16'b0010000001110000: out_v[258] = 10'b1011001010;
    16'b0011000000110000: out_v[258] = 10'b0000111100;
    16'b0010000001010000: out_v[258] = 10'b0110110100;
    16'b0000000000000000: out_v[258] = 10'b0011000100;
    16'b0010000000000000: out_v[258] = 10'b0010110111;
    16'b0010000000110010: out_v[258] = 10'b1111001110;
    16'b0010000001110010: out_v[258] = 10'b1010000111;
    16'b0001000000100000: out_v[258] = 10'b0110000110;
    16'b0001000000110000: out_v[258] = 10'b1111000111;
    16'b0000000000000001: out_v[258] = 10'b1010101100;
    16'b0010010010110000: out_v[258] = 10'b0000011101;
    16'b0000000001010000: out_v[258] = 10'b0011001110;
    16'b0011000000010000: out_v[258] = 10'b0110111011;
    16'b0011000000110001: out_v[258] = 10'b0010101101;
    16'b0000000001010001: out_v[258] = 10'b0001011100;
    16'b0011000000100000: out_v[258] = 10'b0110010111;
    16'b0010000010110000: out_v[258] = 10'b1101111100;
    16'b0010000001010001: out_v[258] = 10'b0100000000;
    16'b0000000001000001: out_v[258] = 10'b1100000101;
    16'b0010000011110000: out_v[258] = 10'b0110001101;
    16'b0010000001010011: out_v[258] = 10'b0011011000;
    16'b0000000000010010: out_v[258] = 10'b0001010101;
    16'b0010000001010010: out_v[258] = 10'b0000111110;
    16'b0000000001110010: out_v[258] = 10'b0101110010;
    16'b0000000000010011: out_v[258] = 10'b1110101110;
    16'b0000010011100010: out_v[258] = 10'b0000110010;
    16'b0000010001110010: out_v[258] = 10'b0101110001;
    16'b0000000001110001: out_v[258] = 10'b0011110010;
    16'b0010000000010010: out_v[258] = 10'b1111001100;
    16'b0000000000110010: out_v[258] = 10'b0001111111;
    16'b0000010010110010: out_v[258] = 10'b1111010001;
    16'b0000000000100000: out_v[258] = 10'b0011110010;
    16'b0010010010010010: out_v[258] = 10'b0111100010;
    16'b0000000001000000: out_v[258] = 10'b1111000101;
    16'b0000000001010010: out_v[258] = 10'b0010011111;
    16'b0000010011010010: out_v[258] = 10'b1001110011;
    16'b0000010011110010: out_v[258] = 10'b0001011001;
    16'b0000000001110011: out_v[258] = 10'b1000011001;
    16'b0000000000100010: out_v[258] = 10'b0000110101;
    16'b0000000000100001: out_v[258] = 10'b0010110100;
    16'b0000000000000010: out_v[258] = 10'b0011010110;
    16'b0000000001100000: out_v[258] = 10'b0100011100;
    16'b0010000010010010: out_v[258] = 10'b1111000111;
    16'b0000000010110010: out_v[258] = 10'b0111110010;
    16'b0000000011110010: out_v[258] = 10'b0000110010;
    16'b0010010011110010: out_v[258] = 10'b1100100000;
    16'b0000000000110011: out_v[258] = 10'b0000111110;
    16'b0010010010110010: out_v[258] = 10'b1111010010;
    16'b0000000001010011: out_v[258] = 10'b0111011001;
    16'b0000000001000010: out_v[258] = 10'b0101011011;
    16'b0000000001110000: out_v[258] = 10'b0011011001;
    16'b0000010010100010: out_v[258] = 10'b0110011101;
    16'b0010000000010011: out_v[258] = 10'b0110101011;
    16'b0000010011000010: out_v[258] = 10'b1100111010;
    16'b0000000000100011: out_v[258] = 10'b0011100000;
    16'b0010000000110011: out_v[258] = 10'b1010001110;
    16'b0010010011010010: out_v[258] = 10'b1000110000;
    16'b0011000000010001: out_v[258] = 10'b0011010011;
    16'b0011000000000001: out_v[258] = 10'b1011000000;
    16'b0011000001000001: out_v[258] = 10'b1001100010;
    16'b0011000001010001: out_v[258] = 10'b1001100001;
    16'b0011000001010011: out_v[258] = 10'b0111001000;
    16'b0000000011010010: out_v[258] = 10'b1100011101;
    16'b0000010010010010: out_v[258] = 10'b1101010010;
    16'b0001000001010000: out_v[258] = 10'b1011110010;
    16'b0011000001000011: out_v[258] = 10'b1101110110;
    16'b0011000001010010: out_v[258] = 10'b1011010111;
    16'b0001000001010010: out_v[258] = 10'b1001011111;
    16'b0000010011100011: out_v[258] = 10'b0110101011;
    16'b0000010011101011: out_v[258] = 10'b0110111110;
    16'b0000010010100001: out_v[258] = 10'b1011101001;
    16'b0000010010000011: out_v[258] = 10'b0010000111;
    16'b0000000000001001: out_v[258] = 10'b1101000011;
    16'b0000010000100011: out_v[258] = 10'b1001100001;
    16'b0000010010000001: out_v[258] = 10'b1001011111;
    16'b0000010011000011: out_v[258] = 10'b1010100001;
    16'b0000010010100011: out_v[258] = 10'b0010111111;
    16'b0000000010000001: out_v[258] = 10'b0010111010;
    16'b0000010010001001: out_v[258] = 10'b1111111010;
    16'b0000000000000011: out_v[258] = 10'b1011001011;
    16'b0000000000001000: out_v[258] = 10'b0111111001;
    16'b0000000010100001: out_v[258] = 10'b1111111000;
    16'b0000000010101001: out_v[258] = 10'b1101111011;
    16'b0000010010100000: out_v[258] = 10'b1011101101;
    16'b0000010011101001: out_v[258] = 10'b1101100000;
    16'b0000010010101001: out_v[258] = 10'b1101111111;
    16'b0000010010101011: out_v[258] = 10'b0110111111;
    16'b0000010011100001: out_v[258] = 10'b1101110010;
    16'b0000010011000001: out_v[258] = 10'b0010101110;
    16'b0000000010110001: out_v[258] = 10'b0011110111;
    16'b0000000011100001: out_v[258] = 10'b1111011000;
    16'b0000010010110001: out_v[258] = 10'b0110011011;
    16'b0000000000101000: out_v[258] = 10'b0111111110;
    16'b0000000000101001: out_v[258] = 10'b0011101100;
    16'b0010010011110011: out_v[258] = 10'b1101100010;
    16'b0010010010110011: out_v[258] = 10'b1101010110;
    16'b0010000010010000: out_v[258] = 10'b0110101011;
    16'b0000000000111010: out_v[258] = 10'b1001001111;
    16'b0010000000000010: out_v[258] = 10'b1101111010;
    16'b0000000000011001: out_v[258] = 10'b1010000101;
    16'b0000000000011000: out_v[258] = 10'b1101101001;
    16'b0000000000111011: out_v[258] = 10'b1100101101;
    16'b0000010011110011: out_v[258] = 10'b1111100010;
    16'b0000000000011010: out_v[258] = 10'b1001100111;
    default: out_v[258] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100000100000010: out_v[259] = 10'b0000011010;
    16'b0000010100000010: out_v[259] = 10'b0000111011;
    16'b0100110100000010: out_v[259] = 10'b1000001001;
    16'b0100010100000000: out_v[259] = 10'b1111010010;
    16'b0000000100000010: out_v[259] = 10'b1000001111;
    16'b0100110100010010: out_v[259] = 10'b1100100001;
    16'b0000010100000000: out_v[259] = 10'b0101010011;
    16'b0100110000000000: out_v[259] = 10'b0100001101;
    16'b0100000100000000: out_v[259] = 10'b0100101000;
    16'b0000010000000000: out_v[259] = 10'b0000010101;
    16'b0000110000000000: out_v[259] = 10'b1010111010;
    16'b0000110100000000: out_v[259] = 10'b1011101011;
    16'b0100110100000000: out_v[259] = 10'b1001100011;
    16'b0100010100000010: out_v[259] = 10'b0010010111;
    16'b0100010000000000: out_v[259] = 10'b1011000110;
    16'b0100100100000000: out_v[259] = 10'b0011100001;
    16'b0100110100010000: out_v[259] = 10'b0001101100;
    16'b0000110100000010: out_v[259] = 10'b1011011000;
    16'b0000000100000000: out_v[259] = 10'b1001100010;
    16'b0100000100010000: out_v[259] = 10'b0010010111;
    16'b0000000000000000: out_v[259] = 10'b0001011011;
    16'b0100100100010000: out_v[259] = 10'b0000101001;
    16'b0100000000000000: out_v[259] = 10'b1010000101;
    16'b0000000000010000: out_v[259] = 10'b0011011101;
    16'b0100100100010010: out_v[259] = 10'b0000010111;
    16'b0000100100100010: out_v[259] = 10'b0110000111;
    16'b0000000100100010: out_v[259] = 10'b1000011001;
    16'b0100000000000010: out_v[259] = 10'b1101000001;
    16'b0000000100110010: out_v[259] = 10'b1111111111;
    16'b0000100100110010: out_v[259] = 10'b0101010100;
    16'b0100100000010000: out_v[259] = 10'b0010000111;
    16'b0100100100000010: out_v[259] = 10'b0110011010;
    16'b0000100100010010: out_v[259] = 10'b1100000110;
    16'b0000010100100010: out_v[259] = 10'b1010100111;
    16'b0100000100010010: out_v[259] = 10'b1011001100;
    16'b0000000000000010: out_v[259] = 10'b0110100000;
    16'b0000000100010010: out_v[259] = 10'b1100010111;
    16'b0000100100000010: out_v[259] = 10'b1110011100;
    16'b0000100000010000: out_v[259] = 10'b0101101101;
    16'b0001000000000010: out_v[259] = 10'b0010001011;
    16'b0100100100110010: out_v[259] = 10'b1110111011;
    16'b0001000100000010: out_v[259] = 10'b0001001101;
    16'b0100100000000000: out_v[259] = 10'b1001000101;
    16'b0000000000100000: out_v[259] = 10'b0001011100;
    16'b0100100000010010: out_v[259] = 10'b0110110101;
    16'b0100100100100010: out_v[259] = 10'b1011100100;
    16'b0100000100100010: out_v[259] = 10'b1010111011;
    16'b0000100000000000: out_v[259] = 10'b1101010010;
    16'b0000100000110000: out_v[259] = 10'b1110110010;
    16'b0000000100100000: out_v[259] = 10'b1110011100;
    16'b0000110000000010: out_v[259] = 10'b0011001010;
    16'b0000110000010000: out_v[259] = 10'b1101011010;
    16'b0100110000000010: out_v[259] = 10'b0001100000;
    16'b0101000100000010: out_v[259] = 10'b1000001111;
    16'b0000100100000000: out_v[259] = 10'b1111110101;
    16'b0100010000000010: out_v[259] = 10'b1101110000;
    16'b0000010000000010: out_v[259] = 10'b0011000100;
    16'b0100110000010000: out_v[259] = 10'b0001011000;
    16'b0100110000100010: out_v[259] = 10'b1110101110;
    16'b0000000000100010: out_v[259] = 10'b1101001001;
    16'b0100100000000010: out_v[259] = 10'b1111000011;
    16'b0000110000100000: out_v[259] = 10'b1010101001;
    16'b0000010000100010: out_v[259] = 10'b1011001011;
    16'b0100110000100000: out_v[259] = 10'b1110010101;
    16'b0100000000100010: out_v[259] = 10'b1111101010;
    16'b0100010000100010: out_v[259] = 10'b0011101110;
    16'b0000010000100000: out_v[259] = 10'b1010011100;
    16'b0100000000100000: out_v[259] = 10'b1011000010;
    16'b0100010000100000: out_v[259] = 10'b1111111111;
    16'b0100100000100000: out_v[259] = 10'b1101110000;
    16'b0100110000110000: out_v[259] = 10'b0011110111;
    16'b0100100000100010: out_v[259] = 10'b1011011000;
    16'b0110000100000110: out_v[259] = 10'b1010010110;
    16'b0110000100000111: out_v[259] = 10'b1001011111;
    default: out_v[259] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001101000000000: out_v[260] = 10'b0100011111;
    16'b0011101000110100: out_v[260] = 10'b0010111001;
    16'b0011101000110101: out_v[260] = 10'b0011001011;
    16'b0011001000110100: out_v[260] = 10'b0000100100;
    16'b0011100000000100: out_v[260] = 10'b1011001011;
    16'b0011101000010100: out_v[260] = 10'b0110110110;
    16'b0010100000000000: out_v[260] = 10'b0010001111;
    16'b0000001000110000: out_v[260] = 10'b0010111100;
    16'b0000001000000000: out_v[260] = 10'b1001100101;
    16'b0011001000110101: out_v[260] = 10'b1000011111;
    16'b0010101000110100: out_v[260] = 10'b1100000111;
    16'b0011000000000100: out_v[260] = 10'b0001111010;
    16'b0001101000110100: out_v[260] = 10'b0101010001;
    16'b0011101000000101: out_v[260] = 10'b1101011111;
    16'b0001001000110100: out_v[260] = 10'b1000100110;
    16'b0011101000000100: out_v[260] = 10'b1001011000;
    16'b0011001000010100: out_v[260] = 10'b1001110111;
    16'b0010100000000100: out_v[260] = 10'b1111011100;
    16'b0001101000110000: out_v[260] = 10'b0011000111;
    16'b0010001000110100: out_v[260] = 10'b1110100001;
    16'b0000101000111000: out_v[260] = 10'b1110100000;
    16'b0011001000000100: out_v[260] = 10'b1110100001;
    16'b0010001000010100: out_v[260] = 10'b1010011110;
    16'b0010101000110000: out_v[260] = 10'b1101011000;
    16'b0000101000000000: out_v[260] = 10'b0101011011;
    16'b0000100000000000: out_v[260] = 10'b0100101100;
    16'b0010101000110101: out_v[260] = 10'b1111011101;
    16'b0011101000000000: out_v[260] = 10'b1111100111;
    16'b0010001000110101: out_v[260] = 10'b0110010111;
    16'b0011001000000000: out_v[260] = 10'b0010100111;
    16'b0010101000010100: out_v[260] = 10'b1111110111;
    16'b0010001000000100: out_v[260] = 10'b1101001101;
    16'b0011100000000101: out_v[260] = 10'b0010001000;
    16'b0010101000000100: out_v[260] = 10'b1110000111;
    16'b0011101000100100: out_v[260] = 10'b0111111000;
    16'b0011101000111100: out_v[260] = 10'b1011101001;
    16'b0001001000000000: out_v[260] = 10'b1000010111;
    16'b0000101000001000: out_v[260] = 10'b1010011111;
    16'b0000100000001000: out_v[260] = 10'b1001101111;
    16'b0000101000110000: out_v[260] = 10'b0001110110;
    16'b0000001000111000: out_v[260] = 10'b1000101010;
    16'b0000000000000000: out_v[260] = 10'b0110101011;
    16'b0000000000001000: out_v[260] = 10'b1010100110;
    16'b0000101000100000: out_v[260] = 10'b0011011101;
    16'b0000101000101000: out_v[260] = 10'b0110100100;
    16'b0000000000111000: out_v[260] = 10'b0000010111;
    16'b0000001000001000: out_v[260] = 10'b0000101100;
    16'b0000001000101000: out_v[260] = 10'b0111110001;
    16'b0010001000001000: out_v[260] = 10'b0110110110;
    16'b0000100000001001: out_v[260] = 10'b0011111101;
    16'b0010000000001000: out_v[260] = 10'b0110111010;
    16'b0011001000111100: out_v[260] = 10'b0110100100;
    16'b0010100000001001: out_v[260] = 10'b1101011000;
    16'b0010100000001000: out_v[260] = 10'b0110000111;
    16'b0000101000001001: out_v[260] = 10'b1101110100;
    16'b0010101000001000: out_v[260] = 10'b0111011011;
    16'b0001001000110000: out_v[260] = 10'b0111011011;
    16'b0000001000001001: out_v[260] = 10'b0111100101;
    16'b0001001000111000: out_v[260] = 10'b1011101000;
    16'b0010001000111000: out_v[260] = 10'b1011000010;
    16'b0010100000000001: out_v[260] = 10'b0000011011;
    16'b0001001000111100: out_v[260] = 10'b1100000110;
    16'b0011001000001000: out_v[260] = 10'b0000110111;
    16'b0011001000111000: out_v[260] = 10'b1110001010;
    16'b0001101000111000: out_v[260] = 10'b1110000110;
    16'b0010101000111000: out_v[260] = 10'b0110100100;
    16'b0000001000111001: out_v[260] = 10'b0010010100;
    16'b0010110000000000: out_v[260] = 10'b0010000100;
    16'b0010101000000000: out_v[260] = 10'b1111100010;
    16'b0010110000001000: out_v[260] = 10'b1001001110;
    16'b0010101000001001: out_v[260] = 10'b0110001111;
    16'b0010001000001001: out_v[260] = 10'b0111100001;
    16'b0010101000001100: out_v[260] = 10'b1011010011;
    16'b0011100000001101: out_v[260] = 10'b1101000100;
    16'b0011101000001100: out_v[260] = 10'b0001001011;
    16'b0011101000001101: out_v[260] = 10'b1011011011;
    16'b0000001000011000: out_v[260] = 10'b1100000011;
    16'b0010001000111001: out_v[260] = 10'b1101100011;
    16'b0011100000001100: out_v[260] = 10'b1100001110;
    16'b0010100000001100: out_v[260] = 10'b0000110100;
    16'b0001100000001100: out_v[260] = 10'b0110001110;
    16'b0000001000111100: out_v[260] = 10'b1110000111;
    16'b0001000000001000: out_v[260] = 10'b0011110001;
    16'b0001000000111000: out_v[260] = 10'b0010111011;
    16'b0000000000111100: out_v[260] = 10'b0100111111;
    16'b0001101000001100: out_v[260] = 10'b0000111111;
    16'b0000000000011000: out_v[260] = 10'b0110011000;
    16'b0001100000001000: out_v[260] = 10'b1100010101;
    16'b0000100000001100: out_v[260] = 10'b1010100101;
    16'b0011000000001100: out_v[260] = 10'b0001110010;
    16'b0001000000001100: out_v[260] = 10'b0011010000;
    16'b0001000000111100: out_v[260] = 10'b0110011000;
    16'b0011000000001101: out_v[260] = 10'b1010011110;
    16'b0010000000111000: out_v[260] = 10'b1101001010;
    16'b0000001000001100: out_v[260] = 10'b1000011110;
    16'b0000000000001100: out_v[260] = 10'b0001111011;
    16'b0000001000101100: out_v[260] = 10'b1011111011;
    16'b0000000000110000: out_v[260] = 10'b1001011110;
    16'b0001001000001100: out_v[260] = 10'b0110100100;
    16'b0000101000001100: out_v[260] = 10'b0001111011;
    16'b0001000000000000: out_v[260] = 10'b1011000010;
    16'b0000100000111000: out_v[260] = 10'b0110000000;
    16'b0011000000111100: out_v[260] = 10'b1000110011;
    16'b0001000000011000: out_v[260] = 10'b0101011111;
    16'b0000100000011000: out_v[260] = 10'b1001100101;
    16'b0010001000101000: out_v[260] = 10'b1001100111;
    16'b0000100000010000: out_v[260] = 10'b1001111010;
    16'b0000001000100000: out_v[260] = 10'b0110110110;
    16'b0000100000110000: out_v[260] = 10'b1100100110;
    16'b0010001000000000: out_v[260] = 10'b0110110111;
    16'b0010001000110000: out_v[260] = 10'b1001100010;
    16'b0011001000100100: out_v[260] = 10'b1010110011;
    16'b0010001000100000: out_v[260] = 10'b1011101000;
    16'b0011000000001000: out_v[260] = 10'b0011011110;
    16'b0010000000001100: out_v[260] = 10'b0011001010;
    16'b0010000000000100: out_v[260] = 10'b1111110100;
    16'b0010101000101000: out_v[260] = 10'b1101010110;
    16'b0011001000001100: out_v[260] = 10'b0111110000;
    16'b0011101000101100: out_v[260] = 10'b1001000010;
    16'b0010000000000000: out_v[260] = 10'b0111010000;
    16'b0011010000001100: out_v[260] = 10'b1111000000;
    16'b0001100000011101: out_v[260] = 10'b0111111110;
    16'b0100100000001001: out_v[260] = 10'b0110001001;
    16'b0001100000000001: out_v[260] = 10'b1001110011;
    16'b0001100000000000: out_v[260] = 10'b0111010010;
    16'b0001100000000100: out_v[260] = 10'b1001101011;
    16'b0100100000001000: out_v[260] = 10'b1101101011;
    16'b0000100000011001: out_v[260] = 10'b0011010010;
    16'b0100100000000001: out_v[260] = 10'b1001011111;
    16'b0001100000000101: out_v[260] = 10'b0010011111;
    16'b0001100000011001: out_v[260] = 10'b1101011111;
    16'b0001100000001101: out_v[260] = 10'b0111001111;
    16'b0001100000001001: out_v[260] = 10'b1101011111;
    16'b0001100000011000: out_v[260] = 10'b1001000101;
    16'b0000100000000001: out_v[260] = 10'b1100110111;
    16'b0101100000000001: out_v[260] = 10'b1110111111;
    16'b0011100000000001: out_v[260] = 10'b1111100011;
    16'b0000101000011000: out_v[260] = 10'b1001101101;
    16'b0001001000001000: out_v[260] = 10'b1110001010;
    16'b0001101000111100: out_v[260] = 10'b1100111001;
    16'b0001101000001000: out_v[260] = 10'b0101111000;
    16'b0011100000001000: out_v[260] = 10'b1000001111;
    16'b0100000000001000: out_v[260] = 10'b1111100111;
    default: out_v[260] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1010101110101011: out_v[261] = 10'b0110010011;
    16'b0010101010101001: out_v[261] = 10'b1011000111;
    16'b0001101010001000: out_v[261] = 10'b1110100111;
    16'b1010001100101011: out_v[261] = 10'b0110110110;
    16'b0011101010101001: out_v[261] = 10'b0110110111;
    16'b0000101010101001: out_v[261] = 10'b0111010001;
    16'b0000101000101001: out_v[261] = 10'b1110011011;
    16'b0110101000001001: out_v[261] = 10'b0011011101;
    16'b0101101010001001: out_v[261] = 10'b1011010111;
    16'b1010101010001001: out_v[261] = 10'b0011000100;
    16'b1010001110001011: out_v[261] = 10'b1110111111;
    16'b1001101010101001: out_v[261] = 10'b1010011010;
    16'b1010101110001011: out_v[261] = 10'b1010111111;
    16'b0001101010001001: out_v[261] = 10'b0010111111;
    16'b0001101010101001: out_v[261] = 10'b1011100111;
    16'b1010101010101001: out_v[261] = 10'b1110110010;
    16'b1010101000101001: out_v[261] = 10'b1110011010;
    16'b1010101100101011: out_v[261] = 10'b1010001111;
    16'b0000101000011000: out_v[261] = 10'b1110011101;
    16'b0000101000001000: out_v[261] = 10'b1100110111;
    16'b0001101010000000: out_v[261] = 10'b1011000011;
    16'b1010001010101001: out_v[261] = 10'b0011011001;
    16'b1000101010101001: out_v[261] = 10'b1010011001;
    16'b1010001100100011: out_v[261] = 10'b1011010111;
    16'b0001101000001000: out_v[261] = 10'b1001000101;
    16'b0110101010001001: out_v[261] = 10'b0110010111;
    16'b0010101010001001: out_v[261] = 10'b1011000010;
    16'b1010001100000011: out_v[261] = 10'b1110101010;
    16'b1011101010001001: out_v[261] = 10'b0111011011;
    16'b1011101010101001: out_v[261] = 10'b0111011000;
    16'b1010001100001011: out_v[261] = 10'b1111111100;
    16'b1010001110100011: out_v[261] = 10'b0111001011;
    16'b0000100000001000: out_v[261] = 10'b0110101101;
    16'b0010101000101001: out_v[261] = 10'b1101001111;
    16'b0001101010100001: out_v[261] = 10'b0111111010;
    16'b0000101010001000: out_v[261] = 10'b0111110010;
    16'b0000000000000000: out_v[261] = 10'b1101000010;
    16'b1000000000000001: out_v[261] = 10'b0011101001;
    16'b0000000000100001: out_v[261] = 10'b1110111010;
    16'b0010000000100001: out_v[261] = 10'b1110010011;
    16'b1010000000100001: out_v[261] = 10'b1011010111;
    16'b1010000000000001: out_v[261] = 10'b0001101110;
    16'b0000000000000001: out_v[261] = 10'b0001100011;
    16'b1000000000000000: out_v[261] = 10'b1110101001;
    16'b1010000000000000: out_v[261] = 10'b1011000011;
    16'b0100000000000000: out_v[261] = 10'b0101111111;
    16'b0000000000100000: out_v[261] = 10'b1111001100;
    16'b0000001000000000: out_v[261] = 10'b0011100011;
    16'b1011000000000001: out_v[261] = 10'b1101100111;
    16'b1011000000100001: out_v[261] = 10'b1010000010;
    16'b1000000000100001: out_v[261] = 10'b1010101011;
    16'b0010000000000001: out_v[261] = 10'b0110000101;
    16'b0000001010000000: out_v[261] = 10'b1110110010;
    16'b1001001110101011: out_v[261] = 10'b0101111011;
    16'b0001001010001000: out_v[261] = 10'b0101100100;
    16'b1010000000100011: out_v[261] = 10'b1011111110;
    16'b1001001000101001: out_v[261] = 10'b1010001110;
    16'b0001001010000000: out_v[261] = 10'b0011101011;
    16'b1011001010100001: out_v[261] = 10'b0011100110;
    16'b1000001000101011: out_v[261] = 10'b1111111011;
    16'b1001001010101011: out_v[261] = 10'b1010100011;
    16'b1001001010101001: out_v[261] = 10'b0111010100;
    16'b1010001000100001: out_v[261] = 10'b1001111101;
    16'b0001001100001000: out_v[261] = 10'b1110000100;
    16'b1001001010001011: out_v[261] = 10'b1011100111;
    16'b1001001010100001: out_v[261] = 10'b0011111010;
    16'b1011001010101001: out_v[261] = 10'b1110111011;
    16'b1010001000101011: out_v[261] = 10'b1011001000;
    16'b1011001010101011: out_v[261] = 10'b1011001100;
    16'b0001001010101001: out_v[261] = 10'b1000011111;
    16'b1001000010101011: out_v[261] = 10'b1100111011;
    16'b1000001100101011: out_v[261] = 10'b1011110011;
    16'b0001001000000000: out_v[261] = 10'b0101000100;
    16'b1010000010100001: out_v[261] = 10'b1010111011;
    16'b0011001010100001: out_v[261] = 10'b0011010110;
    16'b1000001000101001: out_v[261] = 10'b1010110010;
    16'b1001001010001001: out_v[261] = 10'b1101100110;
    16'b1001000010101001: out_v[261] = 10'b0010011101;
    16'b1010001010100001: out_v[261] = 10'b1010110101;
    16'b1010001000100011: out_v[261] = 10'b0110101111;
    16'b1001001000101011: out_v[261] = 10'b0110110011;
    16'b0001001010100001: out_v[261] = 10'b1100110110;
    16'b1011000010100001: out_v[261] = 10'b1001000100;
    16'b0001001010001010: out_v[261] = 10'b1111001111;
    16'b1001001100101011: out_v[261] = 10'b0011101010;
    16'b1010001010100011: out_v[261] = 10'b1110110011;
    16'b1001001110101001: out_v[261] = 10'b1101011001;
    16'b1110000000001001: out_v[261] = 10'b1111110010;
    16'b1011100000001001: out_v[261] = 10'b1001110011;
    16'b1111000000001001: out_v[261] = 10'b1101110001;
    16'b1010100010101001: out_v[261] = 10'b1101000111;
    16'b1001100010101001: out_v[261] = 10'b1010111100;
    16'b1111000010001001: out_v[261] = 10'b0001100001;
    16'b1011000000001001: out_v[261] = 10'b0100011000;
    16'b1010100000101001: out_v[261] = 10'b1010010111;
    16'b0101000000000001: out_v[261] = 10'b0110001011;
    16'b1110100000001001: out_v[261] = 10'b1011010111;
    16'b1001000000101001: out_v[261] = 10'b1000001101;
    16'b1001000000100001: out_v[261] = 10'b0110011000;
    16'b1111100000001001: out_v[261] = 10'b1011011111;
    16'b1001100000101001: out_v[261] = 10'b1110001011;
    16'b1101000000000001: out_v[261] = 10'b0110010011;
    16'b1001100000100001: out_v[261] = 10'b0111000111;
    16'b1011100000101001: out_v[261] = 10'b0001000101;
    16'b1010000010101001: out_v[261] = 10'b0101111010;
    16'b0101000000000000: out_v[261] = 10'b0100011100;
    16'b1011000000101001: out_v[261] = 10'b0111011001;
    16'b1110100010001001: out_v[261] = 10'b1011100110;
    16'b1011100010101001: out_v[261] = 10'b0011001011;
    16'b0011000000001000: out_v[261] = 10'b0000001011;
    16'b1000100010101001: out_v[261] = 10'b1000110100;
    16'b1010100000001001: out_v[261] = 10'b0011111011;
    16'b1111100010001001: out_v[261] = 10'b1111100110;
    16'b1101000000001001: out_v[261] = 10'b0111010011;
    16'b1011000010101001: out_v[261] = 10'b0111101000;
    16'b1011001000101001: out_v[261] = 10'b0010001011;
    16'b1010000000101001: out_v[261] = 10'b1110011110;
    16'b1010000000001001: out_v[261] = 10'b0111011010;
    16'b1001000000000001: out_v[261] = 10'b0100000101;
    16'b0001000010000000: out_v[261] = 10'b1011010010;
    16'b1011101000101001: out_v[261] = 10'b1111001000;
    16'b0011100010000000: out_v[261] = 10'b0011011110;
    16'b0001100000000000: out_v[261] = 10'b1100110100;
    16'b0001000000000000: out_v[261] = 10'b0011000100;
    16'b0001100010000000: out_v[261] = 10'b1001001011;
    16'b0011100000000000: out_v[261] = 10'b1101010110;
    16'b0011000000000000: out_v[261] = 10'b0110100000;
    16'b0001100010000001: out_v[261] = 10'b1010001110;
    16'b0011000010001000: out_v[261] = 10'b0111110011;
    16'b0011000010000000: out_v[261] = 10'b1001000010;
    16'b0000100000000000: out_v[261] = 10'b1010000101;
    16'b0101100010000000: out_v[261] = 10'b1111000110;
    16'b1011100010000000: out_v[261] = 10'b0001111111;
    16'b0011100000000001: out_v[261] = 10'b0011100110;
    16'b0011100010001000: out_v[261] = 10'b1110000000;
    16'b0011100000001000: out_v[261] = 10'b0110100111;
    16'b0001101000000000: out_v[261] = 10'b0101111010;
    16'b0001100010001000: out_v[261] = 10'b1111011010;
    16'b1011100000000000: out_v[261] = 10'b0000011011;
    16'b0100100010000000: out_v[261] = 10'b1001001101;
    16'b0011101010001000: out_v[261] = 10'b1110001010;
    16'b0011001010000000: out_v[261] = 10'b1000111000;
    16'b0011101000000000: out_v[261] = 10'b1010101011;
    16'b1001100010000001: out_v[261] = 10'b1111001111;
    16'b1011100010001000: out_v[261] = 10'b0000110101;
    16'b0001100010010000: out_v[261] = 10'b0100011011;
    16'b0011101010000000: out_v[261] = 10'b0111010110;
    16'b0000100010000000: out_v[261] = 10'b0000110101;
    16'b0001000010001000: out_v[261] = 10'b0001011011;
    16'b1001100010000000: out_v[261] = 10'b0011101111;
    16'b1011101010001000: out_v[261] = 10'b0110110011;
    16'b0011001010001000: out_v[261] = 10'b0011110100;
    16'b0000100000010000: out_v[261] = 10'b1001011010;
    16'b0000101000010000: out_v[261] = 10'b0010111011;
    16'b0001100000011000: out_v[261] = 10'b0111101111;
    16'b0111100000001000: out_v[261] = 10'b1111110011;
    16'b0110100000000000: out_v[261] = 10'b1011011111;
    16'b0010100000000000: out_v[261] = 10'b0011101101;
    16'b0101100000000000: out_v[261] = 10'b0110110110;
    16'b0001100000001000: out_v[261] = 10'b0110100010;
    16'b0100100000010000: out_v[261] = 10'b0001110111;
    16'b0010100000001000: out_v[261] = 10'b0111100110;
    16'b0001001000010000: out_v[261] = 10'b0001100011;
    16'b0011100000001001: out_v[261] = 10'b0000111110;
    16'b0000101000000000: out_v[261] = 10'b0011011010;
    16'b0001101000010000: out_v[261] = 10'b0100101010;
    16'b0111100000000000: out_v[261] = 10'b1101010011;
    16'b0111100000001001: out_v[261] = 10'b1101011001;
    16'b0001100000010000: out_v[261] = 10'b0101001111;
    16'b0100100000000000: out_v[261] = 10'b1001100111;
    16'b0000001000010000: out_v[261] = 10'b0010111001;
    16'b0000000000010000: out_v[261] = 10'b1000100100;
    16'b0011100000101001: out_v[261] = 10'b0111010110;
    16'b0011101000001000: out_v[261] = 10'b0001011011;
    16'b1000101010001001: out_v[261] = 10'b1101011011;
    16'b0001001000001000: out_v[261] = 10'b1000010011;
    16'b0001101000101001: out_v[261] = 10'b1011000110;
    16'b1001101000101001: out_v[261] = 10'b1110110111;
    16'b0011101000101001: out_v[261] = 10'b1111011010;
    16'b1001101110101001: out_v[261] = 10'b1100001010;
    16'b1000101110101011: out_v[261] = 10'b1101011111;
    16'b0001100000101001: out_v[261] = 10'b0110100110;
    16'b1000100000101001: out_v[261] = 10'b1110011110;
    16'b1000100010001000: out_v[261] = 10'b1111001111;
    16'b0000100010101001: out_v[261] = 10'b1111110011;
    16'b0001000000101001: out_v[261] = 10'b1101001101;
    16'b0001000000100001: out_v[261] = 10'b1001001101;
    16'b0001000000100000: out_v[261] = 10'b0011101101;
    16'b0001000000001000: out_v[261] = 10'b0001011011;
    16'b0000100000101001: out_v[261] = 10'b1001011001;
    16'b1000101010001000: out_v[261] = 10'b1011011010;
    16'b0010100000101001: out_v[261] = 10'b1111001011;
    16'b1001101110101011: out_v[261] = 10'b1010111110;
    16'b1001101100101011: out_v[261] = 10'b0110100110;
    16'b0101100010010000: out_v[261] = 10'b1011001111;
    16'b0010100010001000: out_v[261] = 10'b0111101110;
    16'b0101000010000000: out_v[261] = 10'b0000110011;
    16'b0010000010001000: out_v[261] = 10'b1010011000;
    16'b0101000010001000: out_v[261] = 10'b0011100010;
    16'b0000000010000000: out_v[261] = 10'b0110000000;
    16'b0100000010000000: out_v[261] = 10'b0001111011;
    16'b0100101010010000: out_v[261] = 10'b1110101111;
    16'b1011100010001001: out_v[261] = 10'b0110000011;
    16'b1010100010000001: out_v[261] = 10'b1011101011;
    16'b0000101010010000: out_v[261] = 10'b0101001010;
    16'b0010100000000001: out_v[261] = 10'b1111011001;
    16'b0100001010000001: out_v[261] = 10'b1011100101;
    16'b0100101010000001: out_v[261] = 10'b1010111110;
    16'b1010100000000001: out_v[261] = 10'b0100011100;
    16'b0100101010000000: out_v[261] = 10'b0010011011;
    16'b0000001010100001: out_v[261] = 10'b0110101010;
    16'b1011100000000001: out_v[261] = 10'b1011001101;
    16'b1011100010000001: out_v[261] = 10'b1101100010;
    16'b0000001010010000: out_v[261] = 10'b1101011010;
    16'b0010100010000001: out_v[261] = 10'b0110110100;
    16'b0100001010000000: out_v[261] = 10'b0101110101;
    16'b0011100010000001: out_v[261] = 10'b0110111100;
    16'b0100001010010000: out_v[261] = 10'b1100001111;
    16'b0001000011001000: out_v[261] = 10'b1101100101;
    16'b0101101010000000: out_v[261] = 10'b1000001110;
    default: out_v[261] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1000000100100000: out_v[262] = 10'b0101110001;
    16'b1000001000100000: out_v[262] = 10'b1001001111;
    16'b1000000100100010: out_v[262] = 10'b0001111001;
    16'b1000000000000000: out_v[262] = 10'b0101110100;
    16'b1000000100000010: out_v[262] = 10'b1001100110;
    16'b1000100100000000: out_v[262] = 10'b0001100111;
    16'b1000100100000010: out_v[262] = 10'b1010010001;
    16'b1000100000000000: out_v[262] = 10'b1111001011;
    16'b0000100000100010: out_v[262] = 10'b0110010100;
    16'b1000000000100000: out_v[262] = 10'b0111001001;
    16'b1000100000000010: out_v[262] = 10'b0011100011;
    16'b1000101100100010: out_v[262] = 10'b1100010101;
    16'b1000001100100010: out_v[262] = 10'b0010101110;
    16'b1000001100100000: out_v[262] = 10'b0011100101;
    16'b0000000100100010: out_v[262] = 10'b0101000000;
    16'b1000000000100010: out_v[262] = 10'b1010000111;
    16'b1000000100000000: out_v[262] = 10'b1000000010;
    16'b1000000000000010: out_v[262] = 10'b0011000110;
    16'b0000001100100010: out_v[262] = 10'b0001110111;
    16'b0000100100100010: out_v[262] = 10'b1010001011;
    16'b0000000000100010: out_v[262] = 10'b1110110010;
    16'b1000001000000000: out_v[262] = 10'b0110011010;
    16'b0000100100000010: out_v[262] = 10'b1110011011;
    16'b0000101100100010: out_v[262] = 10'b1010110011;
    16'b1000100100100010: out_v[262] = 10'b1010000111;
    16'b0000000000000000: out_v[262] = 10'b1000111001;
    16'b0000000000100000: out_v[262] = 10'b1000000010;
    16'b0000000100000010: out_v[262] = 10'b1001000001;
    16'b1000101100100000: out_v[262] = 10'b1101000011;
    16'b0000100000000010: out_v[262] = 10'b1011110110;
    16'b0000000000000010: out_v[262] = 10'b0011100101;
    16'b0000001000000000: out_v[262] = 10'b1100001010;
    16'b0000000100000000: out_v[262] = 10'b0010100110;
    16'b0000000100100000: out_v[262] = 10'b0010000010;
    16'b0000001000100000: out_v[262] = 10'b0100101010;
    16'b1000000000001010: out_v[262] = 10'b1110100110;
    16'b1000000000001000: out_v[262] = 10'b0001001100;
    16'b1000000000010000: out_v[262] = 10'b1111001110;
    16'b0000000000010000: out_v[262] = 10'b0010110000;
    16'b1000000100010010: out_v[262] = 10'b0011100010;
    16'b1000000000110010: out_v[262] = 10'b1111100011;
    16'b0000000000001000: out_v[262] = 10'b1000001100;
    16'b1000000100001010: out_v[262] = 10'b1000111111;
    16'b0000000000010010: out_v[262] = 10'b0100011011;
    16'b1000000000010010: out_v[262] = 10'b0110010010;
    16'b0000000000110000: out_v[262] = 10'b1100000111;
    16'b0000000000001010: out_v[262] = 10'b0111100101;
    16'b1000000000011010: out_v[262] = 10'b0110100111;
    16'b0000001000100010: out_v[262] = 10'b0100010111;
    16'b0000001100000000: out_v[262] = 10'b0111011001;
    16'b1000001100110000: out_v[262] = 10'b1110110011;
    16'b1000001100110010: out_v[262] = 10'b0001011101;
    16'b1000001000110010: out_v[262] = 10'b0111011111;
    16'b1000001000110000: out_v[262] = 10'b1010100010;
    16'b0000001100100000: out_v[262] = 10'b0011001100;
    16'b0000000000110010: out_v[262] = 10'b0001110010;
    16'b1000001000100010: out_v[262] = 10'b1011000000;
    16'b0000001000110010: out_v[262] = 10'b1110000010;
    16'b0000000100110010: out_v[262] = 10'b0001011110;
    16'b1000000000110000: out_v[262] = 10'b1000000110;
    16'b1000001100000000: out_v[262] = 10'b0111110010;
    16'b0000001100110010: out_v[262] = 10'b1010110101;
    16'b1000000100110010: out_v[262] = 10'b0001111101;
    16'b1000000110000000: out_v[262] = 10'b0010110101;
    16'b1000100000010010: out_v[262] = 10'b0101000110;
    16'b1000000100001000: out_v[262] = 10'b1011001000;
    16'b1000000110000010: out_v[262] = 10'b1111101011;
    16'b1000000010000000: out_v[262] = 10'b1110000111;
    16'b1000100000001010: out_v[262] = 10'b0111110100;
    16'b1000000010000010: out_v[262] = 10'b0010001101;
    16'b0000000100001010: out_v[262] = 10'b0111100011;
    16'b1000000100110000: out_v[262] = 10'b0110010110;
    16'b0000000100010000: out_v[262] = 10'b0000101101;
    16'b0000000100110000: out_v[262] = 10'b1011101011;
    16'b1000000100010000: out_v[262] = 10'b0110110011;
    16'b0000001100110000: out_v[262] = 10'b1111000011;
    16'b0000001100010000: out_v[262] = 10'b0111110000;
    16'b0000101100100000: out_v[262] = 10'b0101101000;
    default: out_v[262] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001000000001011: out_v[263] = 10'b0100100111;
    16'b1010001000001110: out_v[263] = 10'b1110111111;
    16'b1000001000001010: out_v[263] = 10'b1111001001;
    16'b1000000000001010: out_v[263] = 10'b1000001101;
    16'b0000000000001011: out_v[263] = 10'b0110011111;
    16'b1000001000001110: out_v[263] = 10'b0011101111;
    16'b0011001000001011: out_v[263] = 10'b0110110001;
    16'b0000001000000011: out_v[263] = 10'b0101011001;
    16'b1000000000001011: out_v[263] = 10'b0011001100;
    16'b0000001000001011: out_v[263] = 10'b1111010011;
    16'b0011000000001011: out_v[263] = 10'b0011111001;
    16'b1000000000001111: out_v[263] = 10'b0011111110;
    16'b1000000000001110: out_v[263] = 10'b0110100110;
    16'b1000001100001010: out_v[263] = 10'b1001111010;
    16'b1001000000001011: out_v[263] = 10'b1000100011;
    16'b1000000000001001: out_v[263] = 10'b1001010111;
    16'b1000000100001010: out_v[263] = 10'b1011010111;
    16'b0000000000001010: out_v[263] = 10'b1100001101;
    16'b0000001100001110: out_v[263] = 10'b1111001111;
    16'b1000001000001111: out_v[263] = 10'b0111100001;
    16'b0011000000000011: out_v[263] = 10'b1001100101;
    16'b1000000100000110: out_v[263] = 10'b1000011001;
    16'b1000001000001011: out_v[263] = 10'b1001011011;
    16'b1010001000001011: out_v[263] = 10'b0011011110;
    16'b1011000000001011: out_v[263] = 10'b0001101000;
    16'b1000001100001110: out_v[263] = 10'b0101000111;
    16'b0011001000000011: out_v[263] = 10'b0011110110;
    16'b0011000000001001: out_v[263] = 10'b1011001000;
    16'b0011001000000001: out_v[263] = 10'b1111100011;
    16'b1011001000001011: out_v[263] = 10'b1000100011;
    16'b1000000100001110: out_v[263] = 10'b1000000100;
    16'b1000000100000010: out_v[263] = 10'b1001001011;
    16'b1010001000001010: out_v[263] = 10'b1111011111;
    16'b0011000000001010: out_v[263] = 10'b1010100111;
    16'b1010000000001011: out_v[263] = 10'b0101110011;
    16'b0001000000001010: out_v[263] = 10'b0101011001;
    16'b1001000000001010: out_v[263] = 10'b1111100010;
    16'b0011000000000010: out_v[263] = 10'b0010010011;
    16'b1000001100000110: out_v[263] = 10'b1111000101;
    16'b0011000000000001: out_v[263] = 10'b1111001011;
    16'b1000000000001000: out_v[263] = 10'b0000111100;
    16'b1001001000001011: out_v[263] = 10'b0100111010;
    16'b0000001000001010: out_v[263] = 10'b0111010110;
    16'b1000000000000010: out_v[263] = 10'b0011100000;
    16'b0000000100001110: out_v[263] = 10'b1011100011;
    16'b1000001000000011: out_v[263] = 10'b1001010010;
    16'b0011000000000000: out_v[263] = 10'b1011101011;
    16'b0010000000000000: out_v[263] = 10'b0110101111;
    16'b0010000000001010: out_v[263] = 10'b0100110011;
    16'b0010000000000010: out_v[263] = 10'b0100011011;
    16'b0000000000000000: out_v[263] = 10'b1100001010;
    16'b1010000000001010: out_v[263] = 10'b0101010011;
    16'b0010000000001000: out_v[263] = 10'b1110001001;
    16'b1011000000001010: out_v[263] = 10'b1100001100;
    16'b0001000000000000: out_v[263] = 10'b1100111100;
    16'b0011000100001010: out_v[263] = 10'b1110001110;
    16'b0000000100001010: out_v[263] = 10'b1011110100;
    16'b0000000000000001: out_v[263] = 10'b0101010111;
    16'b0000000000000010: out_v[263] = 10'b1011000001;
    16'b0000000000001000: out_v[263] = 10'b1101010110;
    16'b1000000000000011: out_v[263] = 10'b1011000011;
    16'b0000000100000000: out_v[263] = 10'b1111100011;
    16'b0000000000001101: out_v[263] = 10'b0101110110;
    16'b0000000000000011: out_v[263] = 10'b1001000100;
    16'b0000000100000010: out_v[263] = 10'b0010111011;
    16'b1000000000000110: out_v[263] = 10'b0010010110;
    16'b0000000001001011: out_v[263] = 10'b1111010111;
    16'b0001001000000011: out_v[263] = 10'b1110001111;
    16'b0000000100001000: out_v[263] = 10'b1111011101;
    16'b0000000000000111: out_v[263] = 10'b1111110110;
    16'b0000001000000001: out_v[263] = 10'b1111101011;
    16'b0000000000001111: out_v[263] = 10'b0010100110;
    16'b1011000000000111: out_v[263] = 10'b0100001100;
    16'b1000000000000111: out_v[263] = 10'b0111101000;
    16'b0000000100001100: out_v[263] = 10'b0011001011;
    16'b0000000000000100: out_v[263] = 10'b0000011011;
    16'b0000000000000101: out_v[263] = 10'b0001011011;
    16'b0001000000000001: out_v[263] = 10'b0110100111;
    16'b0000000000001110: out_v[263] = 10'b0010101001;
    16'b0001001000000001: out_v[263] = 10'b1000100110;
    16'b0000001000000010: out_v[263] = 10'b0110010011;
    16'b0001000000000011: out_v[263] = 10'b0101011010;
    16'b0000000000001001: out_v[263] = 10'b0110111110;
    16'b0000000100000100: out_v[263] = 10'b1100101101;
    16'b0001000000000010: out_v[263] = 10'b0101011000;
    16'b1011000000001111: out_v[263] = 10'b0101011000;
    16'b0011000100001011: out_v[263] = 10'b0001011001;
    16'b0011000000000111: out_v[263] = 10'b1110110111;
    16'b0011000000001000: out_v[263] = 10'b0011101010;
    16'b0011000100000110: out_v[263] = 10'b0111010111;
    16'b0011000101000010: out_v[263] = 10'b1111111111;
    16'b1011000100000111: out_v[263] = 10'b1001011111;
    16'b0011000101001110: out_v[263] = 10'b1011110000;
    16'b0011000000001110: out_v[263] = 10'b0100010110;
    16'b1011000101001110: out_v[263] = 10'b1011011111;
    16'b0001000000001001: out_v[263] = 10'b0000101011;
    16'b1011000100001111: out_v[263] = 10'b0011001001;
    16'b0011000100000111: out_v[263] = 10'b1010011101;
    16'b1001000000001111: out_v[263] = 10'b1001100011;
    16'b0011000000001111: out_v[263] = 10'b0111110101;
    16'b0011000001001010: out_v[263] = 10'b1110110110;
    16'b0010000000001011: out_v[263] = 10'b0010100101;
    16'b1011000000001110: out_v[263] = 10'b1101001100;
    16'b1011000101001111: out_v[263] = 10'b1110011010;
    16'b1011000100000110: out_v[263] = 10'b1001001100;
    16'b0011000000001100: out_v[263] = 10'b0011011110;
    16'b1011000100001110: out_v[263] = 10'b1100111100;
    16'b0011000101001010: out_v[263] = 10'b1010001011;
    16'b0011000101000110: out_v[263] = 10'b1001110111;
    16'b0010000000001001: out_v[263] = 10'b1010001010;
    16'b1001000000001110: out_v[263] = 10'b1000101000;
    16'b0001000000001000: out_v[263] = 10'b1101001000;
    16'b1001000000000000: out_v[263] = 10'b0001011011;
    16'b0000000100000101: out_v[263] = 10'b0010110010;
    16'b0000001100000101: out_v[263] = 10'b0110111010;
    16'b1000000000000000: out_v[263] = 10'b1000011001;
    16'b1001000000000010: out_v[263] = 10'b1100100111;
    16'b1001000000001000: out_v[263] = 10'b0101010011;
    16'b1000000000001101: out_v[263] = 10'b0101111111;
    16'b0000000000001100: out_v[263] = 10'b1001000011;
    16'b1000000000000001: out_v[263] = 10'b0001110011;
    16'b0001000100000101: out_v[263] = 10'b0110011111;
    16'b1000000100000001: out_v[263] = 10'b0110010000;
    16'b0001000000001100: out_v[263] = 10'b0100110100;
    16'b0000001000000000: out_v[263] = 10'b1011001111;
    16'b1000001000000001: out_v[263] = 10'b1111011000;
    16'b0000000101000101: out_v[263] = 10'b0011011110;
    16'b1001000000001001: out_v[263] = 10'b0101100110;
    16'b1001000000001101: out_v[263] = 10'b1001010000;
    16'b1001000000001100: out_v[263] = 10'b0010111100;
    16'b0001001000000000: out_v[263] = 10'b0001100100;
    16'b0001000000001101: out_v[263] = 10'b0000110101;
    16'b1000001000001001: out_v[263] = 10'b1101101001;
    16'b1000001000001101: out_v[263] = 10'b0111010011;
    16'b1000001000000000: out_v[263] = 10'b0111111011;
    16'b1001000100000010: out_v[263] = 10'b0111010001;
    16'b1001000000000011: out_v[263] = 10'b0100110111;
    16'b1001000100001111: out_v[263] = 10'b0110100011;
    16'b1001000100000110: out_v[263] = 10'b0011111010;
    16'b1001000100001011: out_v[263] = 10'b1010110001;
    16'b1001000100000011: out_v[263] = 10'b0011110110;
    16'b1001000100001110: out_v[263] = 10'b1010110011;
    16'b1001000100000111: out_v[263] = 10'b0001101111;
    16'b1001000100001010: out_v[263] = 10'b1011110101;
    16'b1000000000001100: out_v[263] = 10'b0010100100;
    16'b1011000000001000: out_v[263] = 10'b1101010010;
    16'b1010000000001101: out_v[263] = 10'b1111100000;
    16'b1100000000000100: out_v[263] = 10'b1101101001;
    16'b1100000000001110: out_v[263] = 10'b1101011111;
    16'b1010000000001110: out_v[263] = 10'b1110110010;
    16'b1000000001001110: out_v[263] = 10'b1111110011;
    16'b1110000000001101: out_v[263] = 10'b0100011101;
    16'b1010000000001111: out_v[263] = 10'b0111110011;
    16'b1010000000000000: out_v[263] = 10'b1011100011;
    16'b1100000000001111: out_v[263] = 10'b1111110001;
    16'b1100000000001010: out_v[263] = 10'b0111110111;
    16'b1100000000000110: out_v[263] = 10'b0101111110;
    16'b1000000000000100: out_v[263] = 10'b1011100100;
    16'b1010000000000110: out_v[263] = 10'b0111100001;
    16'b1100000000000010: out_v[263] = 10'b1001100101;
    16'b1100000000001100: out_v[263] = 10'b1010010111;
    16'b1010000000000010: out_v[263] = 10'b1101110100;
    16'b1100000000001101: out_v[263] = 10'b0111101001;
    16'b1000000000000101: out_v[263] = 10'b1011100100;
    16'b0000000000000110: out_v[263] = 10'b1101010111;
    16'b1010000000000100: out_v[263] = 10'b1110000111;
    16'b1001000000000110: out_v[263] = 10'b1011100110;
    16'b0001000100000110: out_v[263] = 10'b0111010001;
    16'b1011000000000011: out_v[263] = 10'b0100101111;
    16'b1011000000000010: out_v[263] = 10'b1110001101;
    16'b0001000100000111: out_v[263] = 10'b0101110010;
    16'b1101000000001010: out_v[263] = 10'b1101100011;
    16'b1000000100000111: out_v[263] = 10'b0110100010;
    16'b0101000000001010: out_v[263] = 10'b1101101011;
    16'b1000001100000111: out_v[263] = 10'b1001000000;
    16'b0101000000000010: out_v[263] = 10'b1101101110;
    16'b0000000100000111: out_v[263] = 10'b1000111011;
    16'b1101000000000010: out_v[263] = 10'b1000001110;
    16'b0100000000001010: out_v[263] = 10'b1101010011;
    16'b1000000100000011: out_v[263] = 10'b1010100100;
    default: out_v[263] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000110001001000: out_v[264] = 10'b1100011011;
    16'b0000110101001000: out_v[264] = 10'b0000011010;
    16'b1000110001001000: out_v[264] = 10'b0100011111;
    16'b0000000101000000: out_v[264] = 10'b1110011111;
    16'b0000000100000000: out_v[264] = 10'b1101000001;
    16'b0000010001001000: out_v[264] = 10'b0110000111;
    16'b1000000001001000: out_v[264] = 10'b0001010001;
    16'b0000110101000000: out_v[264] = 10'b1110010011;
    16'b0000110001011000: out_v[264] = 10'b1011011011;
    16'b1000100001001000: out_v[264] = 10'b1110111111;
    16'b0000100101000000: out_v[264] = 10'b1011111000;
    16'b0000110000001000: out_v[264] = 10'b0000111000;
    16'b0000100001001000: out_v[264] = 10'b0010011011;
    16'b0000110100000000: out_v[264] = 10'b1110110110;
    16'b1000110101001000: out_v[264] = 10'b0111111100;
    16'b0000100101001000: out_v[264] = 10'b1010100111;
    16'b0000110101010000: out_v[264] = 10'b0011100011;
    16'b0000010100000000: out_v[264] = 10'b1110011011;
    16'b0000010101010000: out_v[264] = 10'b1101011011;
    16'b0000110101010001: out_v[264] = 10'b0011100011;
    16'b1010110001001000: out_v[264] = 10'b0010111101;
    16'b0000010101000000: out_v[264] = 10'b0111101001;
    16'b0000110100001000: out_v[264] = 10'b1101111110;
    16'b0000110101011001: out_v[264] = 10'b1011111001;
    16'b0000110101011000: out_v[264] = 10'b1111011011;
    16'b0010110001001000: out_v[264] = 10'b0000101011;
    16'b0000010101001000: out_v[264] = 10'b0010001111;
    16'b0000010101010001: out_v[264] = 10'b1101000111;
    16'b0000010100001000: out_v[264] = 10'b0001001101;
    16'b0010110101001000: out_v[264] = 10'b1010001010;
    16'b0000100000001000: out_v[264] = 10'b0010101011;
    16'b1000111001001000: out_v[264] = 10'b1110100110;
    16'b1000111101001000: out_v[264] = 10'b1011101100;
    16'b0010011000000000: out_v[264] = 10'b0110001011;
    16'b0010001000000000: out_v[264] = 10'b1000111100;
    16'b0010001001000000: out_v[264] = 10'b0100000011;
    16'b0010000000000000: out_v[264] = 10'b1000111011;
    16'b0000000000000000: out_v[264] = 10'b0101000110;
    16'b0000001000000000: out_v[264] = 10'b0101000011;
    16'b0010000001000000: out_v[264] = 10'b1000110111;
    16'b0010010000000000: out_v[264] = 10'b0110010011;
    16'b1010011001000000: out_v[264] = 10'b1000001010;
    16'b1010001000000000: out_v[264] = 10'b0000100111;
    16'b1010001001000000: out_v[264] = 10'b1010111110;
    16'b1010011000000000: out_v[264] = 10'b1101000100;
    16'b0010011001000000: out_v[264] = 10'b0101011001;
    16'b0000010000000000: out_v[264] = 10'b1010010100;
    16'b0000011000000000: out_v[264] = 10'b0111001010;
    16'b0010010001000000: out_v[264] = 10'b1011110100;
    16'b0000001001000000: out_v[264] = 10'b0111001000;
    16'b0000000001000000: out_v[264] = 10'b1111010110;
    16'b0010001000010001: out_v[264] = 10'b1001101100;
    16'b1000001000000000: out_v[264] = 10'b0001111010;
    16'b1000001001010000: out_v[264] = 10'b0111110000;
    16'b0000011001000000: out_v[264] = 10'b0000100001;
    16'b1000011001001000: out_v[264] = 10'b1000111100;
    16'b0010001001010001: out_v[264] = 10'b1010110011;
    16'b1000001001001000: out_v[264] = 10'b1011010100;
    16'b0010000000010001: out_v[264] = 10'b1100010100;
    16'b1000001001010001: out_v[264] = 10'b0011100011;
    16'b1000011001000000: out_v[264] = 10'b1000000111;
    16'b1000001000001000: out_v[264] = 10'b1100011111;
    16'b1000111001000000: out_v[264] = 10'b0110010110;
    16'b1000001001011001: out_v[264] = 10'b0010111111;
    16'b1000111001011001: out_v[264] = 10'b0101011100;
    16'b1000101001000000: out_v[264] = 10'b0101010100;
    16'b1000011101001000: out_v[264] = 10'b0101011110;
    16'b1000001001011000: out_v[264] = 10'b1011001011;
    16'b1000001001000000: out_v[264] = 10'b0101101101;
    16'b0000010001000000: out_v[264] = 10'b0011000100;
    16'b0000011001010001: out_v[264] = 10'b1000111111;
    16'b1000101001001000: out_v[264] = 10'b1111000010;
    16'b1000011001010001: out_v[264] = 10'b1110110111;
    16'b1000011001010000: out_v[264] = 10'b1111100011;
    16'b0010000001010001: out_v[264] = 10'b1101110110;
    16'b1000111001010001: out_v[264] = 10'b1010011000;
    16'b1000111000001000: out_v[264] = 10'b1000101000;
    16'b1010001000010001: out_v[264] = 10'b0010010101;
    16'b1000111001010000: out_v[264] = 10'b0101011111;
    16'b1000001000010001: out_v[264] = 10'b1100101011;
    16'b0000011001001000: out_v[264] = 10'b0110100100;
    16'b1000111001011000: out_v[264] = 10'b1110001111;
    16'b1010001001010001: out_v[264] = 10'b1111000001;
    16'b0010010001001000: out_v[264] = 10'b0110010100;
    16'b1010000001010001: out_v[264] = 10'b1111011110;
    16'b1010010001000000: out_v[264] = 10'b1011011010;
    16'b1000000001010001: out_v[264] = 10'b0101111011;
    16'b0010110001000000: out_v[264] = 10'b1011001010;
    16'b1010110001000000: out_v[264] = 10'b0001110100;
    16'b1010001001011001: out_v[264] = 10'b0010111111;
    16'b1010000001010000: out_v[264] = 10'b1101011111;
    16'b1010000000010001: out_v[264] = 10'b1101010011;
    16'b1010010001001000: out_v[264] = 10'b0101011010;
    16'b1010000001000000: out_v[264] = 10'b0110011000;
    16'b1010010001011000: out_v[264] = 10'b0011110011;
    16'b1010000001011001: out_v[264] = 10'b1000111011;
    16'b0010100000010001: out_v[264] = 10'b0101011010;
    16'b1000010001001000: out_v[264] = 10'b1011101011;
    16'b1010100001000000: out_v[264] = 10'b1011011000;
    16'b0010100001000000: out_v[264] = 10'b0100110010;
    16'b1010000000000000: out_v[264] = 10'b0101011010;
    16'b1010010001010001: out_v[264] = 10'b1110011001;
    16'b1010000001001000: out_v[264] = 10'b0111100000;
    16'b1010110001010001: out_v[264] = 10'b0011111111;
    16'b1000000001000000: out_v[264] = 10'b1000110011;
    16'b1010010001010000: out_v[264] = 10'b1100011111;
    16'b1010011001001000: out_v[264] = 10'b1110001100;
    16'b1010001000011001: out_v[264] = 10'b0010000011;
    16'b1000000000010001: out_v[264] = 10'b1101011110;
    16'b1010000000011001: out_v[264] = 10'b1111001110;
    16'b1000000000000000: out_v[264] = 10'b0111110001;
    16'b1010010001011001: out_v[264] = 10'b0111110011;
    16'b1010100001010001: out_v[264] = 10'b0111111111;
    16'b1000010001000000: out_v[264] = 10'b1010011011;
    16'b0010100001011001: out_v[264] = 10'b0110111000;
    16'b0010100001010001: out_v[264] = 10'b1010100010;
    16'b1010011001010000: out_v[264] = 10'b0011111111;
    16'b1010011001010001: out_v[264] = 10'b1100101111;
    16'b1010011001011001: out_v[264] = 10'b0111011011;
    16'b0010110001010001: out_v[264] = 10'b1111111010;
    16'b1010001001010000: out_v[264] = 10'b0011011001;
    16'b1000011000001000: out_v[264] = 10'b0010111100;
    16'b1010001000001000: out_v[264] = 10'b0111100001;
    16'b1000111100001000: out_v[264] = 10'b0001011111;
    16'b1000101100001000: out_v[264] = 10'b1101111011;
    16'b1000111100011001: out_v[264] = 10'b0110010010;
    16'b1000011100011000: out_v[264] = 10'b0010111101;
    16'b1000011000000000: out_v[264] = 10'b0100011011;
    16'b1000001100001000: out_v[264] = 10'b0101011011;
    16'b1000101100011000: out_v[264] = 10'b1001110111;
    16'b1000001101001000: out_v[264] = 10'b0011011011;
    16'b1000101000011000: out_v[264] = 10'b1100101111;
    16'b1000101000001000: out_v[264] = 10'b1101100010;
    16'b1000101100011001: out_v[264] = 10'b1100101101;
    16'b1000011100001000: out_v[264] = 10'b1010010001;
    16'b1000001000011001: out_v[264] = 10'b0011000110;
    16'b1000010000001000: out_v[264] = 10'b0010100110;
    16'b1000011100011001: out_v[264] = 10'b1100110110;
    16'b1000101101001000: out_v[264] = 10'b0111110100;
    16'b1000001000011000: out_v[264] = 10'b0011111111;
    16'b1000111100011000: out_v[264] = 10'b1011011110;
    16'b1000100100001000: out_v[264] = 10'b0110111000;
    16'b1000101100000000: out_v[264] = 10'b1101010110;
    16'b1000111000011000: out_v[264] = 10'b1010001000;
    16'b0000011000001000: out_v[264] = 10'b1011010101;
    16'b1010001001001000: out_v[264] = 10'b1110010001;
    16'b1010011000001000: out_v[264] = 10'b1001000001;
    16'b1000011000011000: out_v[264] = 10'b1000110111;
    16'b1000000000001000: out_v[264] = 10'b0011000000;
    16'b0000001000001000: out_v[264] = 10'b1001110110;
    16'b1000010000000000: out_v[264] = 10'b0100100011;
    16'b0000000000001000: out_v[264] = 10'b0101111100;
    16'b0000010000001000: out_v[264] = 10'b1100110101;
    16'b0010001000001000: out_v[264] = 10'b0110111111;
    16'b1000010100001000: out_v[264] = 10'b1001100100;
    16'b0000100001000000: out_v[264] = 10'b0000111010;
    16'b0010000000001000: out_v[264] = 10'b1000101100;
    16'b1000000001010000: out_v[264] = 10'b1111110010;
    16'b1010010000000000: out_v[264] = 10'b1010100111;
    16'b1001101100011001: out_v[264] = 10'b1011101110;
    16'b0000000001001000: out_v[264] = 10'b1110010111;
    16'b0000101000001000: out_v[264] = 10'b1011000000;
    16'b0000101001001000: out_v[264] = 10'b1001101111;
    16'b1000101101000000: out_v[264] = 10'b1001010011;
    16'b1000100000001000: out_v[264] = 10'b0001010111;
    16'b0000001001001000: out_v[264] = 10'b1101011001;
    16'b0010100000001000: out_v[264] = 10'b0011010101;
    16'b0010100001001000: out_v[264] = 10'b1011010010;
    16'b0000100000000000: out_v[264] = 10'b1111000111;
    16'b1010001000010000: out_v[264] = 10'b0011101001;
    16'b1000011000000100: out_v[264] = 10'b0110100011;
    16'b1000011100000000: out_v[264] = 10'b1011011010;
    16'b1010011000010001: out_v[264] = 10'b0111100001;
    16'b1000011000010000: out_v[264] = 10'b1001110111;
    16'b1000101000010001: out_v[264] = 10'b0110001111;
    16'b1000101000000100: out_v[264] = 10'b0010101010;
    16'b1000100100000000: out_v[264] = 10'b1101001000;
    16'b1000001000000100: out_v[264] = 10'b0011010011;
    16'b1000111000010100: out_v[264] = 10'b1011100110;
    16'b1010101000010001: out_v[264] = 10'b0101100110;
    16'b1000011000010001: out_v[264] = 10'b1010100011;
    16'b1000101000000000: out_v[264] = 10'b0100000111;
    16'b1000001000010000: out_v[264] = 10'b0111011111;
    16'b0000011000000100: out_v[264] = 10'b0011100011;
    16'b1000011000010101: out_v[264] = 10'b1100110111;
    16'b1010100000000000: out_v[264] = 10'b1101011011;
    16'b1000100000000000: out_v[264] = 10'b1001011011;
    16'b1000111000010001: out_v[264] = 10'b0101101100;
    16'b1000111000010101: out_v[264] = 10'b1010100011;
    16'b1000100000010001: out_v[264] = 10'b1010000110;
    16'b1010101000000000: out_v[264] = 10'b0010110011;
    16'b1000111000000100: out_v[264] = 10'b0001011111;
    16'b1010101000000100: out_v[264] = 10'b1101010110;
    16'b1000111000000000: out_v[264] = 10'b0100011100;
    16'b1000101000010101: out_v[264] = 10'b1110011011;
    16'b0010001001001000: out_v[264] = 10'b0110000111;
    16'b0010011001001000: out_v[264] = 10'b1101101000;
    16'b0000111001000000: out_v[264] = 10'b0110010100;
    16'b1000111100000000: out_v[264] = 10'b1101110111;
    16'b1000011000001100: out_v[264] = 10'b1011000001;
    16'b1000111100001100: out_v[264] = 10'b1001000111;
    16'b1000111000001100: out_v[264] = 10'b1001000100;
    16'b1000110100001000: out_v[264] = 10'b1001001110;
    16'b1000000100001000: out_v[264] = 10'b1100111101;
    16'b1010000000001000: out_v[264] = 10'b1101000110;
    16'b1010001100001000: out_v[264] = 10'b0001110011;
    default: out_v[264] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1101101001000010: out_v[265] = 10'b1100010001;
    16'b1101011001000000: out_v[265] = 10'b1110100100;
    16'b0100011001000011: out_v[265] = 10'b1011011010;
    16'b1100000001000011: out_v[265] = 10'b0110011011;
    16'b0100011001000010: out_v[265] = 10'b0000000111;
    16'b0000001001000011: out_v[265] = 10'b1010100110;
    16'b0100101001000010: out_v[265] = 10'b0000011100;
    16'b1101101001000000: out_v[265] = 10'b0000011011;
    16'b0100001001000011: out_v[265] = 10'b0011101011;
    16'b1101001001000011: out_v[265] = 10'b1001011100;
    16'b0100001001000010: out_v[265] = 10'b1010001111;
    16'b0100001001000000: out_v[265] = 10'b0011000001;
    16'b0101001001000010: out_v[265] = 10'b1100000110;
    16'b1100101001000011: out_v[265] = 10'b0111000101;
    16'b0100000001000011: out_v[265] = 10'b1011101011;
    16'b1101001001000000: out_v[265] = 10'b0011011101;
    16'b0100001001000001: out_v[265] = 10'b1001011001;
    16'b1100001001000011: out_v[265] = 10'b1001110010;
    16'b1101011001000011: out_v[265] = 10'b0110110000;
    16'b1101001001000010: out_v[265] = 10'b0011111100;
    16'b1101011001000010: out_v[265] = 10'b1111110100;
    16'b0100101001000011: out_v[265] = 10'b1001011100;
    16'b1100011001000011: out_v[265] = 10'b1000011010;
    16'b1101011000000000: out_v[265] = 10'b0100100111;
    16'b0100100001000011: out_v[265] = 10'b1000101000;
    16'b1100001001000010: out_v[265] = 10'b0001011010;
    16'b1001011000000000: out_v[265] = 10'b0001001001;
    16'b0000001001000001: out_v[265] = 10'b0000111001;
    16'b1101010001000000: out_v[265] = 10'b0001110001;
    16'b0100000001000010: out_v[265] = 10'b1011001100;
    16'b1001000000000000: out_v[265] = 10'b0010110011;
    16'b1101111001000000: out_v[265] = 10'b0001101011;
    16'b1100011001000010: out_v[265] = 10'b1000011101;
    16'b1101111001000010: out_v[265] = 10'b1011010001;
    16'b1001100000000000: out_v[265] = 10'b1111110001;
    16'b1101101001000011: out_v[265] = 10'b1100010101;
    16'b0000001000000011: out_v[265] = 10'b0010110101;
    16'b0000001001000010: out_v[265] = 10'b1011110101;
    16'b1101000001000000: out_v[265] = 10'b0001001011;
    16'b1100100001000011: out_v[265] = 10'b0011011011;
    16'b0000111000000000: out_v[265] = 10'b1011110111;
    16'b1000101000000000: out_v[265] = 10'b1101100110;
    16'b1100000001000000: out_v[265] = 10'b0110110011;
    16'b1100000000000000: out_v[265] = 10'b1101111111;
    16'b0000101000000000: out_v[265] = 10'b1001110011;
    16'b1100001001000000: out_v[265] = 10'b0100110010;
    16'b1000100000000000: out_v[265] = 10'b1101001100;
    16'b1101000000000000: out_v[265] = 10'b0111111011;
    16'b0000110000000000: out_v[265] = 10'b1000010011;
    16'b1000000001000000: out_v[265] = 10'b1111011101;
    16'b1100101001000000: out_v[265] = 10'b0100110011;
    16'b1000000000000000: out_v[265] = 10'b1101101010;
    16'b1000101001000000: out_v[265] = 10'b1111110001;
    16'b1000110000000000: out_v[265] = 10'b1111011001;
    16'b1101100001000000: out_v[265] = 10'b1001011010;
    16'b1000111000000000: out_v[265] = 10'b1010011110;
    16'b1000001001000000: out_v[265] = 10'b1111000000;
    16'b1000001000000000: out_v[265] = 10'b1100000111;
    16'b0000100000000000: out_v[265] = 10'b0001100010;
    16'b1100100001000000: out_v[265] = 10'b0011111010;
    16'b1001111000000000: out_v[265] = 10'b1011011111;
    16'b0000001000000000: out_v[265] = 10'b1101001111;
    16'b0000000001000000: out_v[265] = 10'b0110010111;
    16'b0100101001000000: out_v[265] = 10'b0011110100;
    16'b1100100001000001: out_v[265] = 10'b0010101100;
    16'b0000100001000000: out_v[265] = 10'b0011110100;
    16'b0100100001000000: out_v[265] = 10'b0010111101;
    16'b1100100000000011: out_v[265] = 10'b1000111001;
    16'b0000100001000001: out_v[265] = 10'b1100110001;
    16'b0000000000000000: out_v[265] = 10'b1100010010;
    16'b0000001001000000: out_v[265] = 10'b0010001101;
    16'b0100110001000000: out_v[265] = 10'b0101110111;
    16'b0000110001000000: out_v[265] = 10'b0011110000;
    16'b1000100001000000: out_v[265] = 10'b0100110101;
    16'b0100000001000000: out_v[265] = 10'b0000101111;
    16'b0000100001000011: out_v[265] = 10'b1001101011;
    16'b0100101001000001: out_v[265] = 10'b0101010111;
    16'b0100100001000001: out_v[265] = 10'b1110001011;
    16'b0000101001000000: out_v[265] = 10'b1011110101;
    16'b0100110001000011: out_v[265] = 10'b1101101001;
    16'b0100010001000000: out_v[265] = 10'b0010111110;
    16'b0000101001000011: out_v[265] = 10'b0111001111;
    16'b0100100001000010: out_v[265] = 10'b1001001111;
    16'b0000010000000000: out_v[265] = 10'b1010010110;
    16'b1100100000000000: out_v[265] = 10'b1000100101;
    16'b0000101001000001: out_v[265] = 10'b1110011010;
    16'b1101100001000001: out_v[265] = 10'b1110100110;
    16'b1000100000000011: out_v[265] = 10'b1000101101;
    16'b1101100001000011: out_v[265] = 10'b1100000101;
    16'b1100110001000000: out_v[265] = 10'b1010101110;
    16'b1100100001000010: out_v[265] = 10'b0110001011;
    16'b0100110001000010: out_v[265] = 10'b1110100101;
    16'b0100111001000011: out_v[265] = 10'b1001000100;
    16'b0100100000000011: out_v[265] = 10'b1011101111;
    16'b1001011001000000: out_v[265] = 10'b1100001110;
    16'b0001001001000000: out_v[265] = 10'b1011100100;
    16'b1101001001000001: out_v[265] = 10'b1101001111;
    16'b1001001001000000: out_v[265] = 10'b0000011010;
    16'b0101011001000000: out_v[265] = 10'b1010111100;
    16'b0101001001000000: out_v[265] = 10'b1001101100;
    16'b1101000001000011: out_v[265] = 10'b1011011001;
    16'b1100001001000001: out_v[265] = 10'b1100011110;
    16'b0101001001000001: out_v[265] = 10'b0001110110;
    16'b0101001001000011: out_v[265] = 10'b1001100110;
    16'b1001000001000000: out_v[265] = 10'b0100011001;
    16'b1101000001000001: out_v[265] = 10'b1001011110;
    16'b1001001001000001: out_v[265] = 10'b1011001100;
    16'b1101011001000001: out_v[265] = 10'b1011011101;
    16'b0100011001000000: out_v[265] = 10'b0011010011;
    16'b1001001000000000: out_v[265] = 10'b1010100100;
    16'b0001011001000000: out_v[265] = 10'b1110111110;
    16'b0101011001000011: out_v[265] = 10'b0101111001;
    16'b1101001000000000: out_v[265] = 10'b0011100001;
    16'b0000100000000011: out_v[265] = 10'b0001010000;
    16'b0000001000000010: out_v[265] = 10'b0100011001;
    16'b0000000000000011: out_v[265] = 10'b0101011001;
    16'b0000011000000010: out_v[265] = 10'b1111100011;
    16'b0000000000000001: out_v[265] = 10'b0001011001;
    16'b0000000000000010: out_v[265] = 10'b0101111000;
    16'b0100000000000010: out_v[265] = 10'b0001011011;
    16'b0000010000000010: out_v[265] = 10'b1011000001;
    16'b0001011000000000: out_v[265] = 10'b0111101101;
    16'b0000010000000011: out_v[265] = 10'b1010000011;
    16'b0000110000000011: out_v[265] = 10'b1010010001;
    16'b0000010000000001: out_v[265] = 10'b1011101011;
    16'b0001000000000000: out_v[265] = 10'b0110110101;
    16'b0000111000000010: out_v[265] = 10'b1111101100;
    16'b0000011000000000: out_v[265] = 10'b1100010100;
    16'b0000110000000010: out_v[265] = 10'b1010111011;
    16'b0000000001000011: out_v[265] = 10'b1110010111;
    16'b0000100000000001: out_v[265] = 10'b0001010011;
    16'b0001000000000010: out_v[265] = 10'b0100111111;
    16'b0001000000000011: out_v[265] = 10'b0010110110;
    16'b0000100000000010: out_v[265] = 10'b0001011011;
    16'b0001001000000010: out_v[265] = 10'b0100110110;
    16'b0000011000000011: out_v[265] = 10'b1001011100;
    16'b0000101000000011: out_v[265] = 10'b1100111000;
    16'b0000101000000010: out_v[265] = 10'b0010011001;
    16'b0100001000000010: out_v[265] = 10'b0101001111;
    16'b1000000000000010: out_v[265] = 10'b0011101111;
    16'b1101001000000010: out_v[265] = 10'b1101100010;
    16'b0101000001000011: out_v[265] = 10'b0110100110;
    16'b1000001000000010: out_v[265] = 10'b1011100001;
    16'b0101011001000010: out_v[265] = 10'b1111010110;
    16'b1001001000000010: out_v[265] = 10'b0010101111;
    16'b1001101000000000: out_v[265] = 10'b1001111000;
    16'b0100001000000011: out_v[265] = 10'b1011100100;
    16'b1101001000000011: out_v[265] = 10'b1001000101;
    16'b1101100001000010: out_v[265] = 10'b1001001000;
    16'b1101110001000000: out_v[265] = 10'b1011011100;
    16'b0101100001000000: out_v[265] = 10'b1001010010;
    16'b0001100000000010: out_v[265] = 10'b1111001011;
    16'b1101110001000010: out_v[265] = 10'b1111010111;
    16'b0101100001000010: out_v[265] = 10'b0110110001;
    16'b0001100000000000: out_v[265] = 10'b0110110100;
    16'b1001100001000000: out_v[265] = 10'b0001111010;
    16'b0000100000100011: out_v[265] = 10'b1101011000;
    16'b1001110000000000: out_v[265] = 10'b1011001010;
    16'b0101100000000000: out_v[265] = 10'b1011001000;
    16'b0100100000000010: out_v[265] = 10'b1100110111;
    16'b1001010000000000: out_v[265] = 10'b0001011000;
    16'b0001100000000011: out_v[265] = 10'b1110001001;
    16'b0101100000000010: out_v[265] = 10'b0111111010;
    16'b1001100000000011: out_v[265] = 10'b1111000110;
    16'b0101000001000000: out_v[265] = 10'b1011001101;
    16'b1001000000000010: out_v[265] = 10'b1011000111;
    16'b1100001000000011: out_v[265] = 10'b1110110101;
    16'b1000000000000011: out_v[265] = 10'b1010100010;
    16'b1000101000000011: out_v[265] = 10'b0011001011;
    16'b1100000000000011: out_v[265] = 10'b1111110001;
    16'b1100101000000011: out_v[265] = 10'b0111001010;
    16'b0100000000000011: out_v[265] = 10'b1111000110;
    16'b1100001000000010: out_v[265] = 10'b1100001111;
    16'b1000001000000011: out_v[265] = 10'b1111100000;
    16'b0100000000000001: out_v[265] = 10'b1110000101;
    16'b1100000000000010: out_v[265] = 10'b1100001000;
    16'b1001001000000011: out_v[265] = 10'b0111100110;
    16'b1001000000000011: out_v[265] = 10'b0111001010;
    16'b0100101000000011: out_v[265] = 10'b1110001010;
    16'b0100001000000001: out_v[265] = 10'b1110100001;
    16'b0101101001000000: out_v[265] = 10'b0101100001;
    16'b0101101001000010: out_v[265] = 10'b0010100111;
    16'b0101111001000000: out_v[265] = 10'b0110110010;
    16'b0100111001000010: out_v[265] = 10'b0111000010;
    16'b0101101001000011: out_v[265] = 10'b0111101010;
    16'b0101111001000011: out_v[265] = 10'b1100110011;
    16'b0101111001000010: out_v[265] = 10'b1111011011;
    16'b0001101001000011: out_v[265] = 10'b0110000110;
    16'b1100101001000010: out_v[265] = 10'b1000111100;
    16'b0101100001000011: out_v[265] = 10'b1110010011;
    16'b1101111001000011: out_v[265] = 10'b1010110001;
    16'b0001101001000010: out_v[265] = 10'b1111101111;
    16'b1100011001000000: out_v[265] = 10'b1111110101;
    16'b1100111001000000: out_v[265] = 10'b0110010001;
    16'b1100100000000010: out_v[265] = 10'b1100001111;
    16'b1100000001000010: out_v[265] = 10'b1101010001;
    16'b0101000001000010: out_v[265] = 10'b0100111001;
    16'b1101000001000010: out_v[265] = 10'b1001100111;
    16'b0100000001000001: out_v[265] = 10'b1111001111;
    16'b1101000000000010: out_v[265] = 10'b0001011001;
    16'b1101000000000011: out_v[265] = 10'b1100011000;
    default: out_v[265] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1000000000010000: out_v[266] = 10'b0101011111;
    16'b0011100000010100: out_v[266] = 10'b0100111110;
    16'b0001100000010100: out_v[266] = 10'b1000011001;
    16'b1000100000010000: out_v[266] = 10'b0101011110;
    16'b0011100000010000: out_v[266] = 10'b1100100011;
    16'b0011000000010100: out_v[266] = 10'b1101010111;
    16'b1010100000010000: out_v[266] = 10'b0100100001;
    16'b1011100000010000: out_v[266] = 10'b0001001110;
    16'b0011000000010000: out_v[266] = 10'b1101010110;
    16'b1011100010010000: out_v[266] = 10'b1011001110;
    16'b0101100000000100: out_v[266] = 10'b1111001110;
    16'b0001000000010000: out_v[266] = 10'b1011100011;
    16'b0111100000010100: out_v[266] = 10'b1101010101;
    16'b0001100000000000: out_v[266] = 10'b0011111011;
    16'b0001100000010000: out_v[266] = 10'b0100000011;
    16'b0001000000000000: out_v[266] = 10'b0101110101;
    16'b0011000000000100: out_v[266] = 10'b0111010011;
    16'b0001100000000100: out_v[266] = 10'b1010010100;
    16'b0111100000000100: out_v[266] = 10'b1011000010;
    16'b0101100000010100: out_v[266] = 10'b0101100111;
    16'b0001000000000100: out_v[266] = 10'b0011001001;
    16'b1011100000010100: out_v[266] = 10'b1110011011;
    16'b1001100010010100: out_v[266] = 10'b0011101001;
    16'b1001100000010100: out_v[266] = 10'b0111001001;
    16'b0101000000000100: out_v[266] = 10'b0101110111;
    16'b0001100010010000: out_v[266] = 10'b1011001111;
    16'b1001100000010000: out_v[266] = 10'b1110100110;
    16'b0011100000000100: out_v[266] = 10'b0111000110;
    16'b0001000000010100: out_v[266] = 10'b0111111001;
    16'b0011100000000000: out_v[266] = 10'b0111001011;
    16'b1011000000010000: out_v[266] = 10'b1010111000;
    16'b1010000000010000: out_v[266] = 10'b0001101011;
    16'b1001100010010000: out_v[266] = 10'b0001010011;
    16'b1011100010010100: out_v[266] = 10'b1001110001;
    16'b0000100000010000: out_v[266] = 10'b0110001011;
    16'b0011100010010000: out_v[266] = 10'b1000101001;
    16'b0111000000000100: out_v[266] = 10'b0101011011;
    16'b1011000010000000: out_v[266] = 10'b1001100101;
    16'b1010000010000000: out_v[266] = 10'b0010101010;
    16'b0000000010000000: out_v[266] = 10'b0011000110;
    16'b1010000000000000: out_v[266] = 10'b0110101100;
    16'b0000000000000000: out_v[266] = 10'b0011011010;
    16'b1011000000000000: out_v[266] = 10'b0010010100;
    16'b1000000010000000: out_v[266] = 10'b0011111101;
    16'b0010000010000000: out_v[266] = 10'b0011101100;
    16'b1000000000000000: out_v[266] = 10'b0011010011;
    16'b0000000010010000: out_v[266] = 10'b1010110101;
    16'b1010000010010000: out_v[266] = 10'b0110011001;
    16'b1000000010010000: out_v[266] = 10'b0101001000;
    16'b0010000010010000: out_v[266] = 10'b1101100100;
    16'b1110000010000001: out_v[266] = 10'b0011111011;
    16'b1111000010000001: out_v[266] = 10'b0010011110;
    16'b0001100010000000: out_v[266] = 10'b0111000110;
    16'b1111000010000000: out_v[266] = 10'b0011100101;
    16'b1011000000000001: out_v[266] = 10'b1100001011;
    16'b0011000010000000: out_v[266] = 10'b1000011011;
    16'b1011000010000001: out_v[266] = 10'b1010100101;
    16'b1110000000000001: out_v[266] = 10'b0110110100;
    16'b1110000000000000: out_v[266] = 10'b1001010110;
    16'b1001000010010000: out_v[266] = 10'b0100100110;
    16'b1001000010000000: out_v[266] = 10'b0100010100;
    16'b0011000010000001: out_v[266] = 10'b1111100101;
    16'b1101100010000000: out_v[266] = 10'b0111101010;
    16'b1011100010000000: out_v[266] = 10'b0110110101;
    16'b1101000010000000: out_v[266] = 10'b0000000101;
    16'b1110000010000000: out_v[266] = 10'b1001111111;
    16'b0111000010000000: out_v[266] = 10'b1011011011;
    16'b1010000010000001: out_v[266] = 10'b1111110000;
    16'b1011000010010000: out_v[266] = 10'b1111011100;
    16'b1111000000000000: out_v[266] = 10'b1011110100;
    16'b0001000010000000: out_v[266] = 10'b0011101010;
    16'b1101000010000001: out_v[266] = 10'b0011111111;
    16'b1001000010000001: out_v[266] = 10'b0101011111;
    16'b1111000010010000: out_v[266] = 10'b1011100110;
    16'b1010100010000000: out_v[266] = 10'b1100100101;
    16'b1111000000000001: out_v[266] = 10'b0111111010;
    16'b0111000010000001: out_v[266] = 10'b1011001101;
    16'b1001100010000000: out_v[266] = 10'b0110010110;
    16'b1001000000000000: out_v[266] = 10'b0101001100;
    16'b1000100010000000: out_v[266] = 10'b0100110001;
    16'b0011000000000000: out_v[266] = 10'b0001011001;
    16'b0100000000010001: out_v[266] = 10'b1111111011;
    16'b0010000000010000: out_v[266] = 10'b1000001110;
    16'b0010000000000000: out_v[266] = 10'b0000011010;
    16'b0000000000010000: out_v[266] = 10'b0100100001;
    16'b0111000000000001: out_v[266] = 10'b1011110111;
    16'b0010000010000001: out_v[266] = 10'b1011110001;
    16'b0111000000000000: out_v[266] = 10'b1011011011;
    16'b0110000010000000: out_v[266] = 10'b0000011111;
    16'b0011000010010000: out_v[266] = 10'b1001100100;
    16'b0010100000010000: out_v[266] = 10'b1111101100;
    16'b0011000000000001: out_v[266] = 10'b0111110100;
    16'b0010000000000001: out_v[266] = 10'b0111010100;
    16'b0011000000010001: out_v[266] = 10'b0101010100;
    16'b0011100000010001: out_v[266] = 10'b0011111110;
    16'b0001000000010001: out_v[266] = 10'b1111011111;
    16'b0111000000010001: out_v[266] = 10'b0011110111;
    16'b0000000000010001: out_v[266] = 10'b1011011001;
    16'b0010100000000000: out_v[266] = 10'b1011110111;
    16'b0011100010000000: out_v[266] = 10'b1010101111;
    16'b0101000000010001: out_v[266] = 10'b0011110101;
    16'b0110000000000000: out_v[266] = 10'b0011001111;
    16'b0110000010000001: out_v[266] = 10'b0101011101;
    16'b0010100010000000: out_v[266] = 10'b1000000101;
    16'b1010100010010000: out_v[266] = 10'b1100111010;
    16'b0010100010010000: out_v[266] = 10'b0011111111;
    16'b0000100010010000: out_v[266] = 10'b0010011001;
    16'b0110100010000001: out_v[266] = 10'b1011001111;
    16'b0000100010000000: out_v[266] = 10'b1011010011;
    16'b0010100010010100: out_v[266] = 10'b0100011010;
    16'b0110100000000000: out_v[266] = 10'b1111100011;
    16'b0110100010000000: out_v[266] = 10'b1101000001;
    16'b0000100000000000: out_v[266] = 10'b1001110000;
    16'b1000100010010000: out_v[266] = 10'b1100001110;
    16'b0100100010000000: out_v[266] = 10'b1101100000;
    16'b1110100010000000: out_v[266] = 10'b1111101010;
    16'b1010100010010100: out_v[266] = 10'b0000110011;
    16'b0010100010000100: out_v[266] = 10'b1000010111;
    16'b1110100010000001: out_v[266] = 10'b0100101011;
    16'b0001000010010000: out_v[266] = 10'b1010101010;
    16'b0101000000010000: out_v[266] = 10'b0010110001;
    16'b0101100000010000: out_v[266] = 10'b1011100111;
    16'b0100100000000000: out_v[266] = 10'b1001100111;
    16'b0101100000000000: out_v[266] = 10'b0111000110;
    16'b1001000000010000: out_v[266] = 10'b0110100100;
    16'b1000100010000101: out_v[266] = 10'b1111101010;
    16'b1000100010010100: out_v[266] = 10'b0100110001;
    16'b1000100010000100: out_v[266] = 10'b0101001110;
    16'b1000000010010100: out_v[266] = 10'b1010101110;
    16'b0001100010010100: out_v[266] = 10'b1011111111;
    16'b1100100010010000: out_v[266] = 10'b0011110110;
    16'b1000100000000100: out_v[266] = 10'b1111001011;
    16'b1000100000010100: out_v[266] = 10'b1000000011;
    16'b1010100010000100: out_v[266] = 10'b1010111110;
    16'b1000100000000000: out_v[266] = 10'b0110111010;
    16'b0010000100010000: out_v[266] = 10'b1111010111;
    16'b0010000110010000: out_v[266] = 10'b1011010110;
    16'b1110000010010000: out_v[266] = 10'b0011100101;
    16'b1110000000010000: out_v[266] = 10'b1011101001;
    16'b1110100010010000: out_v[266] = 10'b1110110111;
    default: out_v[266] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0011001110000100: out_v[267] = 10'b0010000101;
    16'b0010001100000000: out_v[267] = 10'b0110110011;
    16'b0001000100000100: out_v[267] = 10'b0100111011;
    16'b1000000110000100: out_v[267] = 10'b0101100011;
    16'b0001000110000100: out_v[267] = 10'b1110110111;
    16'b0010000100000000: out_v[267] = 10'b0011110001;
    16'b0000000010000100: out_v[267] = 10'b0000000011;
    16'b0000000000000100: out_v[267] = 10'b0010110011;
    16'b0011000100000100: out_v[267] = 10'b1100011110;
    16'b1001000000000100: out_v[267] = 10'b1111100111;
    16'b0011011100000000: out_v[267] = 10'b1001000111;
    16'b0000000000000000: out_v[267] = 10'b0110011011;
    16'b0000000110000100: out_v[267] = 10'b0011111000;
    16'b0010000100000100: out_v[267] = 10'b0011001011;
    16'b0000000100000100: out_v[267] = 10'b0010100111;
    16'b0010000110000100: out_v[267] = 10'b0111110111;
    16'b0000000010000000: out_v[267] = 10'b0110100111;
    16'b1011000100000100: out_v[267] = 10'b1100110011;
    16'b0010000010000100: out_v[267] = 10'b1101010110;
    16'b0010001100000100: out_v[267] = 10'b1001001110;
    16'b1001000110000100: out_v[267] = 10'b0110001101;
    16'b0001000000000100: out_v[267] = 10'b0010100001;
    16'b0001000010000100: out_v[267] = 10'b1001000111;
    16'b0000000100000000: out_v[267] = 10'b0011110010;
    16'b0011001000000000: out_v[267] = 10'b0110010011;
    16'b0000001000000100: out_v[267] = 10'b1000001011;
    16'b0011001100000100: out_v[267] = 10'b0000111011;
    16'b0011001100000000: out_v[267] = 10'b0010010011;
    16'b0000001000000000: out_v[267] = 10'b1110100100;
    16'b1000000010000100: out_v[267] = 10'b0111011111;
    16'b0010001000000000: out_v[267] = 10'b1001100011;
    16'b0010001110000100: out_v[267] = 10'b1101110110;
    16'b0000001010000100: out_v[267] = 10'b1010001101;
    16'b1000000000000100: out_v[267] = 10'b1110001001;
    16'b1001000100000100: out_v[267] = 10'b0111000011;
    16'b0011000110000100: out_v[267] = 10'b0100010100;
    16'b0001001000000100: out_v[267] = 10'b0000011101;
    16'b1011000000000100: out_v[267] = 10'b1000001101;
    16'b0000001110000100: out_v[267] = 10'b0100110110;
    16'b0000001100000100: out_v[267] = 10'b0001101110;
    16'b1000000100000100: out_v[267] = 10'b0001100101;
    16'b0001001110000100: out_v[267] = 10'b1011000011;
    16'b0010000000000100: out_v[267] = 10'b0110011101;
    16'b0000001100000000: out_v[267] = 10'b0011100011;
    16'b0001011100000000: out_v[267] = 10'b1111001010;
    16'b0001010100000000: out_v[267] = 10'b1101011110;
    16'b0000010000000000: out_v[267] = 10'b1001001110;
    16'b0000010010000000: out_v[267] = 10'b0111110011;
    16'b0000011000000000: out_v[267] = 10'b1001000101;
    16'b0001010000000000: out_v[267] = 10'b1001100110;
    16'b0001011000000000: out_v[267] = 10'b1000101011;
    16'b0000011010000000: out_v[267] = 10'b0001001101;
    16'b0000011010000100: out_v[267] = 10'b1110100000;
    16'b0001001000000000: out_v[267] = 10'b1111001000;
    16'b0000001010000000: out_v[267] = 10'b1011001011;
    16'b0001010010000000: out_v[267] = 10'b0010110101;
    16'b0011000100000000: out_v[267] = 10'b0011011110;
    16'b0011010100000000: out_v[267] = 10'b0101100000;
    16'b0001010000000100: out_v[267] = 10'b0011111111;
    16'b0011010000000000: out_v[267] = 10'b1100011000;
    16'b0011010110000000: out_v[267] = 10'b1011110111;
    16'b1011011100000000: out_v[267] = 10'b0011001110;
    16'b0011010110000001: out_v[267] = 10'b1101111001;
    16'b0001011010000000: out_v[267] = 10'b1110110011;
    16'b0011011110000100: out_v[267] = 10'b0110011010;
    16'b0011010110000100: out_v[267] = 10'b0011101101;
    16'b0001010100000100: out_v[267] = 10'b0111000100;
    16'b0001010010000100: out_v[267] = 10'b0011110101;
    16'b0001010000000001: out_v[267] = 10'b0111001100;
    16'b0011000110000000: out_v[267] = 10'b0000011110;
    16'b0011011110000000: out_v[267] = 10'b0010001010;
    16'b0001010110000000: out_v[267] = 10'b0011110101;
    16'b0011010110000101: out_v[267] = 10'b1010000101;
    16'b0011000110000101: out_v[267] = 10'b0111001110;
    16'b0001010110000100: out_v[267] = 10'b0101110001;
    16'b1011010100000000: out_v[267] = 10'b0110001101;
    16'b0001010010000001: out_v[267] = 10'b1110011100;
    16'b0001010110000001: out_v[267] = 10'b0100011010;
    16'b0001011010000100: out_v[267] = 10'b1110000111;
    16'b1011000100000000: out_v[267] = 10'b1011011111;
    16'b0010000110000000: out_v[267] = 10'b0010000110;
    16'b0011010010000000: out_v[267] = 10'b1100100100;
    16'b0001011010000001: out_v[267] = 10'b1010101000;
    16'b0001010010000101: out_v[267] = 10'b0001011110;
    16'b0001011110000000: out_v[267] = 10'b1101010100;
    16'b0011010100000100: out_v[267] = 10'b1010001010;
    16'b0001010110000101: out_v[267] = 10'b1011111111;
    16'b0010011010000100: out_v[267] = 10'b1010010111;
    16'b0010011000000000: out_v[267] = 10'b0001111000;
    16'b0010011010000000: out_v[267] = 10'b0001001110;
    16'b0000011110000000: out_v[267] = 10'b0111001011;
    16'b0010010110000000: out_v[267] = 10'b1111011010;
    16'b0010011100000000: out_v[267] = 10'b0100010100;
    16'b0010011110000000: out_v[267] = 10'b1000011010;
    16'b0010011000000100: out_v[267] = 10'b0010101110;
    16'b0011011010000000: out_v[267] = 10'b1010111010;
    16'b0010011110000100: out_v[267] = 10'b1110010110;
    16'b0010001110000000: out_v[267] = 10'b0100001111;
    16'b0010010010000000: out_v[267] = 10'b1111001001;
    16'b0011011000000000: out_v[267] = 10'b0111100001;
    16'b0010011100000100: out_v[267] = 10'b1110001110;
    16'b0010011000100000: out_v[267] = 10'b1111001001;
    16'b0000011100000000: out_v[267] = 10'b0101010000;
    16'b0010011010100000: out_v[267] = 10'b0100110111;
    16'b0010011010000010: out_v[267] = 10'b1001100011;
    16'b0011011010000100: out_v[267] = 10'b0101100010;
    16'b0010001010000000: out_v[267] = 10'b1100001111;
    16'b0010010110000100: out_v[267] = 10'b1000111010;
    16'b0000011110000100: out_v[267] = 10'b0101011010;
    16'b0000001110000000: out_v[267] = 10'b0010111110;
    16'b0010000000000000: out_v[267] = 10'b1011010100;
    16'b0011011010100000: out_v[267] = 10'b1010111010;
    16'b0010010000000110: out_v[267] = 10'b0111010000;
    16'b0010010000000100: out_v[267] = 10'b0110001010;
    16'b0011011100000100: out_v[267] = 10'b1101011000;
    16'b0010010100000100: out_v[267] = 10'b1001101101;
    16'b0010011000000010: out_v[267] = 10'b0001010111;
    16'b0000010000000100: out_v[267] = 10'b0111010011;
    16'b0010010000000000: out_v[267] = 10'b1111001001;
    16'b0011010000000100: out_v[267] = 10'b0011001101;
    16'b0010011100000110: out_v[267] = 10'b1101011011;
    16'b1010010100000100: out_v[267] = 10'b1010101011;
    16'b0010010100000110: out_v[267] = 10'b0111011011;
    16'b0010011100000010: out_v[267] = 10'b0010011101;
    16'b0010010010000100: out_v[267] = 10'b0001110011;
    16'b0000011000000100: out_v[267] = 10'b0001110001;
    16'b0010000100000010: out_v[267] = 10'b0101011111;
    16'b0010010100000010: out_v[267] = 10'b1011010111;
    16'b0010010100000000: out_v[267] = 10'b1101101010;
    16'b0000011100000100: out_v[267] = 10'b1100011011;
    16'b1010011100000100: out_v[267] = 10'b0111011011;
    16'b0000010100000100: out_v[267] = 10'b1111001010;
    16'b0011011000000100: out_v[267] = 10'b0100101110;
    16'b0010001000000100: out_v[267] = 10'b1001001100;
    16'b0010011010000110: out_v[267] = 10'b1000000110;
    16'b0010001010000100: out_v[267] = 10'b0011110010;
    16'b0001001100000000: out_v[267] = 10'b0001101010;
    16'b0001011000000100: out_v[267] = 10'b1100011100;
    16'b0011000010000100: out_v[267] = 10'b0101100110;
    16'b0011010010000100: out_v[267] = 10'b1100010011;
    16'b0011000000000100: out_v[267] = 10'b0101100110;
    16'b0001011110000100: out_v[267] = 10'b0101100010;
    16'b0011000000000000: out_v[267] = 10'b0111111011;
    16'b0001011100000100: out_v[267] = 10'b1101001101;
    16'b0011001010000100: out_v[267] = 10'b0011110010;
    16'b0011001000000100: out_v[267] = 10'b1111011110;
    16'b0010000100000110: out_v[267] = 10'b0111010111;
    16'b0000010100000000: out_v[267] = 10'b1101001010;
    16'b0000010010000100: out_v[267] = 10'b1001100001;
    16'b1010000100000100: out_v[267] = 10'b1111011110;
    16'b0001011110000110: out_v[267] = 10'b0110010011;
    16'b0011011110000110: out_v[267] = 10'b0111011000;
    16'b0010010010000110: out_v[267] = 10'b1011001100;
    16'b0010010110000110: out_v[267] = 10'b1111100111;
    16'b0011000110000110: out_v[267] = 10'b1011101010;
    16'b0010011000000110: out_v[267] = 10'b0001100011;
    16'b0010000110000110: out_v[267] = 10'b1101101100;
    default: out_v[267] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000101101100000: out_v[268] = 10'b1111101110;
    16'b0001100001100000: out_v[268] = 10'b1000010100;
    16'b0001000001100000: out_v[268] = 10'b0101010011;
    16'b0000100001100000: out_v[268] = 10'b1010010000;
    16'b0000001111100000: out_v[268] = 10'b0111001110;
    16'b0000101111100000: out_v[268] = 10'b1010100001;
    16'b0001100001000000: out_v[268] = 10'b1111110011;
    16'b0001100000000000: out_v[268] = 10'b0011101011;
    16'b0001001001000000: out_v[268] = 10'b1000100001;
    16'b0000001101100000: out_v[268] = 10'b1011001101;
    16'b0000001111000000: out_v[268] = 10'b0110110110;
    16'b0000100000100000: out_v[268] = 10'b1011101011;
    16'b0001101001100000: out_v[268] = 10'b0100000111;
    16'b0000001011100000: out_v[268] = 10'b1010010100;
    16'b0001001011100000: out_v[268] = 10'b1011010101;
    16'b0001001001100000: out_v[268] = 10'b0000011111;
    16'b0001101011100000: out_v[268] = 10'b1011000110;
    16'b0001001111100000: out_v[268] = 10'b1010011111;
    16'b0001100000100000: out_v[268] = 10'b0101000011;
    16'b0000100101100000: out_v[268] = 10'b1010101111;
    16'b0001100100100000: out_v[268] = 10'b0110110000;
    16'b0000001101000000: out_v[268] = 10'b1001001101;
    16'b0000001110000000: out_v[268] = 10'b0001101100;
    16'b0000101001100000: out_v[268] = 10'b0101110111;
    16'b0001101111100000: out_v[268] = 10'b1001011011;
    16'b0000001001100000: out_v[268] = 10'b0010000111;
    16'b0000100000000000: out_v[268] = 10'b0010101101;
    16'b0001100101100000: out_v[268] = 10'b0011111010;
    16'b0001001011000000: out_v[268] = 10'b0110010100;
    16'b0001000001000000: out_v[268] = 10'b0111100011;
    16'b0000000001100000: out_v[268] = 10'b1010001111;
    16'b0001000101100000: out_v[268] = 10'b1001101101;
    16'b0001001101100000: out_v[268] = 10'b1100011110;
    16'b0001101101100000: out_v[268] = 10'b1111001110;
    16'b0001001111000000: out_v[268] = 10'b1000111100;
    16'b0000100100100000: out_v[268] = 10'b1101110100;
    16'b0001000000000000: out_v[268] = 10'b0011010101;
    16'b0000101011100000: out_v[268] = 10'b1101100001;
    16'b0000000110000000: out_v[268] = 10'b1010100111;
    16'b0000000101100000: out_v[268] = 10'b0011110011;
    16'b0001001101000000: out_v[268] = 10'b0000101010;
    16'b0000000000000000: out_v[268] = 10'b0010100110;
    16'b0000000010000000: out_v[268] = 10'b1100001111;
    16'b0000000100000000: out_v[268] = 10'b0000110010;
    16'b0001000110000000: out_v[268] = 10'b1100011010;
    16'b0001000010000000: out_v[268] = 10'b0110000100;
    16'b0001001110000000: out_v[268] = 10'b0010101011;
    16'b0001001010000000: out_v[268] = 10'b1000101100;
    16'b0001000010100000: out_v[268] = 10'b0110011110;
    16'b0000001010000000: out_v[268] = 10'b0100011101;
    16'b0001000011000000: out_v[268] = 10'b0111000101;
    16'b0000001011000000: out_v[268] = 10'b0010010110;
    16'b0000000001000000: out_v[268] = 10'b0111111000;
    16'b0000000011000000: out_v[268] = 10'b0101011100;
    16'b0001100011000000: out_v[268] = 10'b1000111011;
    16'b0001101011000000: out_v[268] = 10'b1101011110;
    16'b0001001010100000: out_v[268] = 10'b1111001010;
    16'b0000001001000000: out_v[268] = 10'b1110110101;
    16'b0001000100000000: out_v[268] = 10'b0011010110;
    16'b0001000011100000: out_v[268] = 10'b1101001101;
    16'b0001101111000000: out_v[268] = 10'b1000000100;
    16'b0000001010100000: out_v[268] = 10'b1100111100;
    16'b0001000101000000: out_v[268] = 10'b1111000010;
    16'b0001001000000000: out_v[268] = 10'b1111101010;
    16'b0001000001010000: out_v[268] = 10'b0001101010;
    16'b0001100100110000: out_v[268] = 10'b1101001001;
    16'b0000000101000000: out_v[268] = 10'b1101101011;
    16'b0001001100000000: out_v[268] = 10'b1100100000;
    16'b0001100100000000: out_v[268] = 10'b1111001001;
    16'b0001000101010000: out_v[268] = 10'b0101011010;
    16'b0001100101000000: out_v[268] = 10'b0100000110;
    16'b0000001100000000: out_v[268] = 10'b0111101001;
    16'b0000001000000000: out_v[268] = 10'b1101011000;
    16'b0000101011000000: out_v[268] = 10'b0010010010;
    16'b0000100010000000: out_v[268] = 10'b0011011110;
    16'b0000000010100000: out_v[268] = 10'b1001010000;
    16'b0000000110100000: out_v[268] = 10'b0110110011;
    16'b0000100011000000: out_v[268] = 10'b0111101011;
    16'b0000000111000000: out_v[268] = 10'b0010110100;
    16'b0000100111000000: out_v[268] = 10'b1110111010;
    16'b0000100010100000: out_v[268] = 10'b1011111111;
    16'b0000001111000100: out_v[268] = 10'b1110101111;
    16'b0101100010100000: out_v[268] = 10'b0011101111;
    16'b0000000101000100: out_v[268] = 10'b1011001011;
    16'b0101101111100000: out_v[268] = 10'b0101110100;
    16'b0101000001000000: out_v[268] = 10'b1101011011;
    16'b0101101011100000: out_v[268] = 10'b0000010101;
    16'b0101000011000000: out_v[268] = 10'b0101101011;
    16'b0000000110000100: out_v[268] = 10'b0001011000;
    16'b0101001011000000: out_v[268] = 10'b1111001010;
    16'b0000101111100100: out_v[268] = 10'b1001101010;
    16'b0101100001100000: out_v[268] = 10'b1100111011;
    16'b0101001111000000: out_v[268] = 10'b1000011010;
    16'b0000001110000100: out_v[268] = 10'b1101011100;
    16'b0101100000100000: out_v[268] = 10'b1111100111;
    16'b0001100010100000: out_v[268] = 10'b0010110111;
    16'b0101001011100000: out_v[268] = 10'b0101100110;
    16'b0001100011100000: out_v[268] = 10'b1110010110;
    16'b0101100011100000: out_v[268] = 10'b1110111010;
    16'b0000001101000100: out_v[268] = 10'b1100011111;
    16'b0000001110100000: out_v[268] = 10'b1101011111;
    16'b0000001111110000: out_v[268] = 10'b1001110010;
    16'b0000001010010000: out_v[268] = 10'b1100111100;
    16'b0000001111010000: out_v[268] = 10'b1001001100;
    16'b0000001110010000: out_v[268] = 10'b1101111111;
    16'b0000001011110000: out_v[268] = 10'b1011111011;
    16'b0000001011010000: out_v[268] = 10'b0001010001;
    16'b0000000010010000: out_v[268] = 10'b1010000010;
    16'b0000001001010000: out_v[268] = 10'b1101110111;
    16'b0001000110100000: out_v[268] = 10'b0110110000;
    16'b0001000000100000: out_v[268] = 10'b1110000011;
    16'b0000000100100000: out_v[268] = 10'b0110000010;
    16'b0001001110100000: out_v[268] = 10'b0110010000;
    default: out_v[268] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000010000001: out_v[269] = 10'b0100000111;
    16'b1000000111000001: out_v[269] = 10'b0111010101;
    16'b1000001110000001: out_v[269] = 10'b0001001001;
    16'b0000000010000000: out_v[269] = 10'b0101101000;
    16'b0000000110000001: out_v[269] = 10'b0100111000;
    16'b0000000100000001: out_v[269] = 10'b1000111100;
    16'b1000001100000001: out_v[269] = 10'b0100010111;
    16'b1000001111000000: out_v[269] = 10'b0101101111;
    16'b1000001010000000: out_v[269] = 10'b0001101011;
    16'b1000000111000000: out_v[269] = 10'b1010111101;
    16'b1000001110000000: out_v[269] = 10'b0011111000;
    16'b1000001111000001: out_v[269] = 10'b1010110011;
    16'b1000000110000000: out_v[269] = 10'b0111001010;
    16'b1000000010000000: out_v[269] = 10'b0011000001;
    16'b1000000010000001: out_v[269] = 10'b0100011011;
    16'b0000000111000000: out_v[269] = 10'b1011000001;
    16'b0000000110000000: out_v[269] = 10'b1000100110;
    16'b0000000101000000: out_v[269] = 10'b1110100101;
    16'b1000001010000001: out_v[269] = 10'b1010111011;
    16'b1000001000000001: out_v[269] = 10'b1110111001;
    16'b0000000111000001: out_v[269] = 10'b1011111010;
    16'b1000001011000000: out_v[269] = 10'b1000110010;
    16'b1000000110000001: out_v[269] = 10'b0000111111;
    16'b1000000101000001: out_v[269] = 10'b1110101011;
    16'b1000000100000001: out_v[269] = 10'b1101010110;
    16'b0000000100000000: out_v[269] = 10'b1001010110;
    16'b1000000101000000: out_v[269] = 10'b1011001110;
    16'b0000000101000001: out_v[269] = 10'b0111011101;
    16'b1000001000100001: out_v[269] = 10'b1111000111;
    16'b1000001010100001: out_v[269] = 10'b0101011011;
    16'b1000001100000000: out_v[269] = 10'b0001101111;
    16'b0000000001000001: out_v[269] = 10'b0000101010;
    16'b0000000000000001: out_v[269] = 10'b0010110000;
    16'b0000000000000000: out_v[269] = 10'b1010110010;
    16'b0000000110100000: out_v[269] = 10'b0110110111;
    16'b0000000110001001: out_v[269] = 10'b1001111101;
    16'b0000000100001001: out_v[269] = 10'b0001110011;
    16'b0000000011000001: out_v[269] = 10'b0101000100;
    16'b0000100100000001: out_v[269] = 10'b0000000110;
    16'b0000000100001000: out_v[269] = 10'b0010011101;
    16'b0000000110100001: out_v[269] = 10'b0010011100;
    16'b0000000000100001: out_v[269] = 10'b0101001111;
    16'b0000000000100000: out_v[269] = 10'b0010111001;
    16'b0000000010100001: out_v[269] = 10'b0010111111;
    16'b0000000100000101: out_v[269] = 10'b0011001010;
    16'b0000000010000101: out_v[269] = 10'b1011000010;
    16'b0000000111000101: out_v[269] = 10'b1111010101;
    16'b0000000010100000: out_v[269] = 10'b1010000100;
    16'b0000000110000101: out_v[269] = 10'b0011011011;
    16'b1000000000000000: out_v[269] = 10'b0010110110;
    16'b1000000000000001: out_v[269] = 10'b1110011010;
    16'b1000001000000000: out_v[269] = 10'b0111001100;
    16'b1000000100000000: out_v[269] = 10'b1110000010;
    16'b0000000011000000: out_v[269] = 10'b0100100000;
    16'b0000000001100000: out_v[269] = 10'b0101100000;
    16'b1000000011000000: out_v[269] = 10'b0100100111;
    16'b1000100110000000: out_v[269] = 10'b1110111101;
    16'b0000100110000000: out_v[269] = 10'b1000001011;
    16'b1000101100000000: out_v[269] = 10'b1011111011;
    16'b1000101110000000: out_v[269] = 10'b0100111111;
    16'b1000100100000000: out_v[269] = 10'b0111000110;
    16'b0000100100000000: out_v[269] = 10'b1111001010;
    16'b0000100010000000: out_v[269] = 10'b0111110011;
    16'b0001000100000001: out_v[269] = 10'b0010001110;
    16'b0010000010000001: out_v[269] = 10'b1000000111;
    16'b0010000110000001: out_v[269] = 10'b1000001010;
    16'b0010000000100001: out_v[269] = 10'b0011101110;
    16'b0010000110100001: out_v[269] = 10'b1010101011;
    16'b0001000000000001: out_v[269] = 10'b1101001101;
    16'b0001000110000001: out_v[269] = 10'b1100111110;
    16'b0010000010100001: out_v[269] = 10'b1100100110;
    16'b0000000001000000: out_v[269] = 10'b1111100101;
    16'b0000000100100001: out_v[269] = 10'b0101011011;
    default: out_v[269] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000001000000000: out_v[270] = 10'b1010101000;
    16'b1010001000000001: out_v[270] = 10'b1000100001;
    16'b1010001001000000: out_v[270] = 10'b0111000110;
    16'b1010000000000000: out_v[270] = 10'b1111001100;
    16'b0010000001000000: out_v[270] = 10'b1010100011;
    16'b1010000000000001: out_v[270] = 10'b0000100011;
    16'b0010000000000000: out_v[270] = 10'b1011100100;
    16'b1000001000000000: out_v[270] = 10'b0010101100;
    16'b0000000000000000: out_v[270] = 10'b1111000011;
    16'b0010001000000000: out_v[270] = 10'b0100000101;
    16'b1010001000000000: out_v[270] = 10'b0111011011;
    16'b1000000000000000: out_v[270] = 10'b0100011111;
    16'b0010001001000000: out_v[270] = 10'b0100000110;
    16'b1010000001000000: out_v[270] = 10'b0000010011;
    16'b1000001001000000: out_v[270] = 10'b0000111101;
    16'b1000001000000001: out_v[270] = 10'b1010100001;
    16'b0000001001000000: out_v[270] = 10'b1001100101;
    16'b1000000000000001: out_v[270] = 10'b1000100001;
    16'b0000000001000000: out_v[270] = 10'b0101101011;
    16'b1010001001000001: out_v[270] = 10'b1001010000;
    16'b0000000000001000: out_v[270] = 10'b1101000100;
    16'b0000000001001000: out_v[270] = 10'b0000110101;
    16'b0000001000001000: out_v[270] = 10'b0101001001;
    16'b0010000001001000: out_v[270] = 10'b0001101010;
    16'b0010000000001000: out_v[270] = 10'b0001011101;
    16'b1010000000000010: out_v[270] = 10'b0010001110;
    16'b1010000001000010: out_v[270] = 10'b1010010000;
    16'b0010001001001000: out_v[270] = 10'b1110111011;
    16'b0010001000001000: out_v[270] = 10'b1110010111;
    16'b0000001001001000: out_v[270] = 10'b1101111011;
    16'b1000000001000000: out_v[270] = 10'b1100110010;
    16'b1000000000000010: out_v[270] = 10'b0110011101;
    16'b1000001000000010: out_v[270] = 10'b0001011100;
    16'b0000000000000001: out_v[270] = 10'b0000111000;
    16'b0000001000000001: out_v[270] = 10'b0100010101;
    16'b0010000000000001: out_v[270] = 10'b0010011011;
    16'b0010001000000001: out_v[270] = 10'b0101011000;
    16'b1000001001000001: out_v[270] = 10'b1111100010;
    16'b0000000010000000: out_v[270] = 10'b1010101110;
    16'b0010000010000000: out_v[270] = 10'b0100100100;
    16'b0000100000000000: out_v[270] = 10'b1010001011;
    16'b0010001010000000: out_v[270] = 10'b1110110110;
    16'b1010001010000000: out_v[270] = 10'b0110011010;
    default: out_v[270] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010000000000010: out_v[271] = 10'b0101111011;
    16'b0000000000000000: out_v[271] = 10'b1000000111;
    16'b0000000100000000: out_v[271] = 10'b1010010111;
    16'b0010000000000000: out_v[271] = 10'b1101001000;
    16'b0010000000001010: out_v[271] = 10'b1000010110;
    16'b0000000000000010: out_v[271] = 10'b0001101000;
    16'b0000000000001000: out_v[271] = 10'b1101110110;
    16'b0010000000001000: out_v[271] = 10'b0111010100;
    16'b0000000000001010: out_v[271] = 10'b1101000011;
    16'b0000000100001000: out_v[271] = 10'b0101011110;
    16'b0010000100001010: out_v[271] = 10'b1010010100;
    16'b0000000100001010: out_v[271] = 10'b0110011011;
    16'b1010000100001010: out_v[271] = 10'b0111110010;
    16'b0010000100000010: out_v[271] = 10'b1000101100;
    16'b0010010000001010: out_v[271] = 10'b0000110110;
    16'b1010000000001010: out_v[271] = 10'b0011010111;
    16'b1000000100001000: out_v[271] = 10'b1010110100;
    16'b1000000000001000: out_v[271] = 10'b1001011011;
    16'b0010000100000000: out_v[271] = 10'b1001001011;
    16'b0000000100001100: out_v[271] = 10'b1000101001;
    16'b0010000100001000: out_v[271] = 10'b1111000010;
    16'b1010000100000010: out_v[271] = 10'b0010111111;
    16'b1010000100001000: out_v[271] = 10'b0101011110;
    16'b0000000000001100: out_v[271] = 10'b0011110001;
    16'b1010000000000000: out_v[271] = 10'b1110011011;
    16'b1010000000000010: out_v[271] = 10'b1100001110;
    16'b0010000000001110: out_v[271] = 10'b1000100110;
    16'b0110000000001010: out_v[271] = 10'b0000010000;
    16'b0010000000101010: out_v[271] = 10'b0010010110;
    16'b0100000000000000: out_v[271] = 10'b1000111011;
    16'b0100000000001000: out_v[271] = 10'b0001100010;
    16'b0000000000101000: out_v[271] = 10'b1000110000;
    16'b0000000000000100: out_v[271] = 10'b0001110011;
    16'b0000000000100000: out_v[271] = 10'b1010100100;
    16'b0000010000001000: out_v[271] = 10'b0001100001;
    16'b0000010000000000: out_v[271] = 10'b1101010010;
    16'b0010010000001000: out_v[271] = 10'b0011010000;
    16'b0010010000000010: out_v[271] = 10'b0011100000;
    16'b0011000000001110: out_v[271] = 10'b1101001011;
    16'b0010000100011010: out_v[271] = 10'b0111110011;
    16'b0011000100001110: out_v[271] = 10'b0011011100;
    16'b1010000100001110: out_v[271] = 10'b1111010011;
    16'b0010000100001110: out_v[271] = 10'b1011001111;
    16'b0011000000001010: out_v[271] = 10'b1000000111;
    16'b0001000000001110: out_v[271] = 10'b1100101011;
    16'b0011000100001010: out_v[271] = 10'b0110111001;
    16'b0010000000000110: out_v[271] = 10'b0111101011;
    16'b0001000000001100: out_v[271] = 10'b0111000101;
    16'b0000000000001110: out_v[271] = 10'b1101011110;
    16'b0010000000001100: out_v[271] = 10'b1101010110;
    default: out_v[271] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001010011010001: out_v[272] = 10'b0110001001;
    16'b0001010001010001: out_v[272] = 10'b0011010001;
    16'b0001010000010011: out_v[272] = 10'b0011011011;
    16'b0001010001000001: out_v[272] = 10'b0000001101;
    16'b0000010000000000: out_v[272] = 10'b1001010100;
    16'b0001010000010000: out_v[272] = 10'b0110010011;
    16'b0000000000010010: out_v[272] = 10'b1100000011;
    16'b0001010001000011: out_v[272] = 10'b0000100011;
    16'b0001010011000011: out_v[272] = 10'b0110000011;
    16'b0001010000000000: out_v[272] = 10'b0100001111;
    16'b0001000001010001: out_v[272] = 10'b0101111100;
    16'b0001010001010011: out_v[272] = 10'b0000100111;
    16'b0001010011000001: out_v[272] = 10'b1000101100;
    16'b0001010010000000: out_v[272] = 10'b0001011101;
    16'b0001010010000001: out_v[272] = 10'b0011101110;
    16'b0000010001000001: out_v[272] = 10'b1110011011;
    16'b0001000000010000: out_v[272] = 10'b1000100011;
    16'b0001010000000001: out_v[272] = 10'b1101100010;
    16'b0000010001010001: out_v[272] = 10'b0111010101;
    16'b0001010010010000: out_v[272] = 10'b1000110111;
    16'b0001010000000011: out_v[272] = 10'b1111110100;
    16'b0001010010000010: out_v[272] = 10'b0010011001;
    16'b0001010010010011: out_v[272] = 10'b1111001111;
    16'b0001010000010010: out_v[272] = 10'b1101011011;
    16'b0001010000010001: out_v[272] = 10'b0110100100;
    16'b0001000000010011: out_v[272] = 10'b0111011111;
    16'b0001000000010001: out_v[272] = 10'b0101110000;
    16'b0001010010010001: out_v[272] = 10'b0001110111;
    16'b0001010011010011: out_v[272] = 10'b0111011101;
    16'b0000010010010000: out_v[272] = 10'b0100001001;
    16'b0000000000010000: out_v[272] = 10'b0011101111;
    16'b0000010010000000: out_v[272] = 10'b1001100101;
    16'b0000010000010000: out_v[272] = 10'b0011011010;
    16'b0001010000000010: out_v[272] = 10'b0100010110;
    16'b0001010010000011: out_v[272] = 10'b1011101001;
    16'b0001010001010000: out_v[272] = 10'b1011001011;
    16'b0101010001010001: out_v[272] = 10'b0110010010;
    16'b0101000001000001: out_v[272] = 10'b1001000111;
    16'b0101010001000001: out_v[272] = 10'b1001101010;
    16'b0100010000000000: out_v[272] = 10'b0101111001;
    16'b0100010000010000: out_v[272] = 10'b0010000010;
    16'b0100000000010000: out_v[272] = 10'b0010110111;
    16'b0001000001000000: out_v[272] = 10'b1011111111;
    16'b0001000001000001: out_v[272] = 10'b0100111011;
    16'b0100000010010000: out_v[272] = 10'b1010000011;
    16'b0100000000000000: out_v[272] = 10'b0010010101;
    16'b0000010001000000: out_v[272] = 10'b1010100001;
    16'b0101000000000001: out_v[272] = 10'b1000110110;
    16'b0001000000000001: out_v[272] = 10'b1010101000;
    16'b0101010000010000: out_v[272] = 10'b1010001100;
    16'b0000000000000000: out_v[272] = 10'b1101100010;
    16'b0101010001000000: out_v[272] = 10'b1010101111;
    16'b0100010001000000: out_v[272] = 10'b0101001010;
    16'b0001010001000000: out_v[272] = 10'b1001101101;
    16'b0101000001000000: out_v[272] = 10'b1100100101;
    16'b0100010010010000: out_v[272] = 10'b0010001010;
    16'b0000000010010000: out_v[272] = 10'b0110011010;
    16'b0101010000000000: out_v[272] = 10'b1000000100;
    16'b0000000001000000: out_v[272] = 10'b0101100110;
    16'b0101010001010000: out_v[272] = 10'b0010111010;
    16'b0100010010000000: out_v[272] = 10'b0111001000;
    16'b0101010010000000: out_v[272] = 10'b1111101010;
    16'b0101000000000000: out_v[272] = 10'b1000000101;
    16'b0000000001000001: out_v[272] = 10'b0100011101;
    16'b0101000011000001: out_v[272] = 10'b1011000101;
    16'b0001000000000000: out_v[272] = 10'b1111100011;
    16'b0111000000000000: out_v[272] = 10'b0011111001;
    16'b0101010011000001: out_v[272] = 10'b1010101001;
    16'b0100000001000001: out_v[272] = 10'b1110000100;
    16'b0110000000000000: out_v[272] = 10'b1001100101;
    16'b0101000001010001: out_v[272] = 10'b1001100101;
    16'b0101010000000001: out_v[272] = 10'b1000010011;
    16'b0001000011000001: out_v[272] = 10'b0101010000;
    16'b0101010010010000: out_v[272] = 10'b0111011000;
    16'b0100000010000000: out_v[272] = 10'b0110111000;
    16'b0000000010000000: out_v[272] = 10'b0101001000;
    16'b0101010010000001: out_v[272] = 10'b1011101000;
    16'b0101000010000000: out_v[272] = 10'b1001011111;
    16'b0101010011010001: out_v[272] = 10'b0101111010;
    16'b0101010000010001: out_v[272] = 10'b1010011000;
    16'b0100010000000001: out_v[272] = 10'b0101011111;
    16'b0101000011000000: out_v[272] = 10'b0101100011;
    16'b0001000010000000: out_v[272] = 10'b1011110110;
    16'b0100000010000001: out_v[272] = 10'b0011110011;
    16'b0000000000000001: out_v[272] = 10'b1000010010;
    16'b0001000010000001: out_v[272] = 10'b0110110000;
    16'b0100010000010001: out_v[272] = 10'b1010111101;
    16'b0101000010000001: out_v[272] = 10'b1110011101;
    16'b0100000000000001: out_v[272] = 10'b0011110011;
    16'b0001000011000000: out_v[272] = 10'b0111110111;
    16'b0101000000010001: out_v[272] = 10'b1011000001;
    16'b0101000000010000: out_v[272] = 10'b1101101011;
    16'b0000010001010000: out_v[272] = 10'b1010100100;
    16'b0101010010010001: out_v[272] = 10'b0110110110;
    16'b0000010011000001: out_v[272] = 10'b1011111110;
    16'b0000010011000000: out_v[272] = 10'b0010100110;
    16'b0100010011000001: out_v[272] = 10'b0111010010;
    16'b0000000000000010: out_v[272] = 10'b1011000011;
    16'b0100010001010000: out_v[272] = 10'b1110100100;
    16'b0000000000100000: out_v[272] = 10'b1111001000;
    16'b0000000001010000: out_v[272] = 10'b1111010010;
    16'b0100000001000000: out_v[272] = 10'b0011010100;
    16'b0100000000000010: out_v[272] = 10'b0011111110;
    16'b0100000001010000: out_v[272] = 10'b1010111001;
    16'b0100000000100000: out_v[272] = 10'b0111101011;
    16'b0100010001010001: out_v[272] = 10'b1110000001;
    16'b1000000010010000: out_v[272] = 10'b1111000000;
    16'b1000000110010000: out_v[272] = 10'b1001111000;
    16'b0000000110010000: out_v[272] = 10'b0111100011;
    16'b1101010000000000: out_v[272] = 10'b0101001011;
    16'b1100010000010000: out_v[272] = 10'b1010000011;
    16'b1001010000000000: out_v[272] = 10'b1101001110;
    16'b1000010000010000: out_v[272] = 10'b1101110101;
    16'b0000000110000000: out_v[272] = 10'b1110101011;
    16'b1001010000010000: out_v[272] = 10'b1111110110;
    16'b1000010000000000: out_v[272] = 10'b0010001011;
    16'b0001000110000000: out_v[272] = 10'b1011101110;
    16'b1000000000000000: out_v[272] = 10'b1010101010;
    16'b1101010000010000: out_v[272] = 10'b1111110110;
    16'b1000000000010000: out_v[272] = 10'b0110011111;
    16'b0100010001000001: out_v[272] = 10'b1111000010;
    16'b0101010011000000: out_v[272] = 10'b1100100111;
    16'b0101000110000000: out_v[272] = 10'b1000001111;
    16'b0100000110000000: out_v[272] = 10'b1000001011;
    16'b0100000100000000: out_v[272] = 10'b1100001011;
    default: out_v[272] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001011000000000: out_v[273] = 10'b1011001001;
    16'b0001011000100010: out_v[273] = 10'b0111100001;
    16'b0000001000000000: out_v[273] = 10'b0001110101;
    16'b0001011000100000: out_v[273] = 10'b0010001011;
    16'b0001010000000000: out_v[273] = 10'b1001101100;
    16'b0001011000000010: out_v[273] = 10'b1000101001;
    16'b0000001000000010: out_v[273] = 10'b0101010101;
    16'b0001010000000010: out_v[273] = 10'b1100000110;
    16'b0000011000100000: out_v[273] = 10'b1110011000;
    16'b0001010000100000: out_v[273] = 10'b1000101010;
    16'b0000011000000000: out_v[273] = 10'b1110100001;
    16'b0000011000000010: out_v[273] = 10'b1100101000;
    16'b0000011000100010: out_v[273] = 10'b0111111011;
    16'b0001010000100010: out_v[273] = 10'b0110110100;
    16'b0000010000100010: out_v[273] = 10'b0100010011;
    16'b0001001000000000: out_v[273] = 10'b0100011110;
    16'b0000000000100000: out_v[273] = 10'b1111100001;
    16'b0000010000100000: out_v[273] = 10'b0100011011;
    16'b0000010000000000: out_v[273] = 10'b1111100101;
    16'b0000000000100010: out_v[273] = 10'b1001000011;
    16'b0001001000100000: out_v[273] = 10'b1101100011;
    16'b0000000000000000: out_v[273] = 10'b0011010110;
    16'b0000000000000010: out_v[273] = 10'b0000010010;
    16'b0001000000100000: out_v[273] = 10'b1010100100;
    16'b0001000000000000: out_v[273] = 10'b0111011011;
    16'b0000001000100000: out_v[273] = 10'b1111101000;
    16'b0000010000000010: out_v[273] = 10'b1010101100;
    16'b0000001000100010: out_v[273] = 10'b1111001010;
    16'b0010011000100000: out_v[273] = 10'b1100011010;
    16'b0011011000100000: out_v[273] = 10'b0001011111;
    16'b0000100000000000: out_v[273] = 10'b0111010111;
    16'b0001000000000010: out_v[273] = 10'b0100011011;
    16'b0001001000000010: out_v[273] = 10'b0001011011;
    16'b0010000000000000: out_v[273] = 10'b0111010010;
    16'b0100000000000000: out_v[273] = 10'b0111100101;
    16'b0011100000100000: out_v[273] = 10'b0011010001;
    16'b0010001000100000: out_v[273] = 10'b0011001110;
    16'b0011011000000000: out_v[273] = 10'b0011110110;
    16'b0000100000100000: out_v[273] = 10'b0111100110;
    16'b0011001000100000: out_v[273] = 10'b0110111001;
    16'b0010000000100000: out_v[273] = 10'b1010001000;
    16'b0010100000100000: out_v[273] = 10'b0011000111;
    16'b0011000000100000: out_v[273] = 10'b1101001111;
    16'b0000110000100000: out_v[273] = 10'b0101011100;
    16'b0000110000000000: out_v[273] = 10'b1100101111;
    16'b0001110000000000: out_v[273] = 10'b1011000110;
    16'b0001110000100000: out_v[273] = 10'b1001101001;
    16'b0001100000100000: out_v[273] = 10'b1101001010;
    default: out_v[273] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1000000000101000: out_v[274] = 10'b1100100011;
    16'b1000000000000000: out_v[274] = 10'b0001011010;
    16'b1000000000100010: out_v[274] = 10'b0111100000;
    16'b1000010000110010: out_v[274] = 10'b1111010011;
    16'b0000000000000000: out_v[274] = 10'b0010100100;
    16'b0000010000100010: out_v[274] = 10'b1100010011;
    16'b1000000000110010: out_v[274] = 10'b0111110010;
    16'b0000000000000010: out_v[274] = 10'b1011001001;
    16'b1000000000100000: out_v[274] = 10'b1111100011;
    16'b0000000000100010: out_v[274] = 10'b0011001111;
    16'b0000010000100000: out_v[274] = 10'b1110000110;
    16'b1000000000001000: out_v[274] = 10'b0011011010;
    16'b1000000000010000: out_v[274] = 10'b1010101110;
    16'b1000000000101010: out_v[274] = 10'b0011011001;
    16'b1000000000110000: out_v[274] = 10'b1010100011;
    16'b1000000000000010: out_v[274] = 10'b1100100101;
    16'b0000000000100000: out_v[274] = 10'b1001011000;
    16'b0000000000010000: out_v[274] = 10'b0100011111;
    16'b0000000000110000: out_v[274] = 10'b1100110011;
    16'b1000010000100010: out_v[274] = 10'b0011000001;
    16'b0000000000001000: out_v[274] = 10'b0010110110;
    16'b0000000000011000: out_v[274] = 10'b0101001100;
    16'b1000010000000010: out_v[274] = 10'b0111010101;
    16'b0000010000000000: out_v[274] = 10'b0100101001;
    16'b0001000000010000: out_v[274] = 10'b1010000011;
    16'b0001000000011000: out_v[274] = 10'b1001100111;
    16'b0001000000001000: out_v[274] = 10'b0111011010;
    16'b0000000000101010: out_v[274] = 10'b0110010101;
    16'b1000000000011000: out_v[274] = 10'b1011011110;
    16'b0000000000101000: out_v[274] = 10'b0100111100;
    16'b0000010000011000: out_v[274] = 10'b1010110110;
    16'b0000010000001000: out_v[274] = 10'b1110001110;
    16'b1000001000001000: out_v[274] = 10'b1010100110;
    16'b0000000000001010: out_v[274] = 10'b0101010000;
    16'b0000000000111000: out_v[274] = 10'b0110111100;
    16'b0000001000001000: out_v[274] = 10'b0010001110;
    16'b1001000000000000: out_v[274] = 10'b0000001100;
    16'b0001000000000000: out_v[274] = 10'b1110001000;
    16'b0100000000000000: out_v[274] = 10'b0101011101;
    16'b1100000000001000: out_v[274] = 10'b0001111101;
    16'b1100000000000000: out_v[274] = 10'b0000011111;
    16'b1001000000001000: out_v[274] = 10'b0011001011;
    16'b1000001000000000: out_v[274] = 10'b1000011010;
    16'b1000010000000000: out_v[274] = 10'b0111001011;
    16'b1000000000001010: out_v[274] = 10'b1101010000;
    16'b1001000000010000: out_v[274] = 10'b0011100111;
    16'b0100000000001000: out_v[274] = 10'b0000111011;
    16'b0100000000101010: out_v[274] = 10'b1001101011;
    16'b0100000000101000: out_v[274] = 10'b1110110011;
    16'b1000000000111000: out_v[274] = 10'b0111000010;
    16'b0100000000001010: out_v[274] = 10'b0110010000;
    16'b0100000000000010: out_v[274] = 10'b1101110001;
    16'b0000000000011010: out_v[274] = 10'b0100110011;
    16'b1000010000101010: out_v[274] = 10'b1001110011;
    16'b1100000000000010: out_v[274] = 10'b1101110110;
    16'b1000000000010010: out_v[274] = 10'b1110100011;
    16'b1000000010100010: out_v[274] = 10'b1011110100;
    16'b1010000000100000: out_v[274] = 10'b0111100011;
    16'b1010000010100010: out_v[274] = 10'b0001110011;
    16'b1010000000100010: out_v[274] = 10'b0111011110;
    16'b1010000000000000: out_v[274] = 10'b1101011011;
    16'b0000000010100010: out_v[274] = 10'b0011001100;
    16'b1000000000100110: out_v[274] = 10'b0111111111;
    16'b1010000000000010: out_v[274] = 10'b0010011111;
    16'b0100000010100010: out_v[274] = 10'b0011101111;
    16'b0010000000100010: out_v[274] = 10'b1011000111;
    16'b1100000000101000: out_v[274] = 10'b0011110100;
    16'b1100000000001010: out_v[274] = 10'b0100010010;
    16'b1100000000101010: out_v[274] = 10'b1100100011;
    16'b1010000000101000: out_v[274] = 10'b1100110111;
    16'b1010000000101010: out_v[274] = 10'b1011011111;
    16'b0010000000101010: out_v[274] = 10'b1001111111;
    16'b0010000000101000: out_v[274] = 10'b0110101111;
    default: out_v[274] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100000000000010: out_v[275] = 10'b1101001000;
    16'b1100000000010001: out_v[275] = 10'b1110001111;
    16'b1100000000000001: out_v[275] = 10'b1100011111;
    16'b1100000000000011: out_v[275] = 10'b1000011011;
    16'b1100000000000010: out_v[275] = 10'b0000011010;
    16'b0100000010000001: out_v[275] = 10'b0000111010;
    16'b0100000010010001: out_v[275] = 10'b1000110101;
    16'b1000000000000011: out_v[275] = 10'b0011111000;
    16'b0100000010000011: out_v[275] = 10'b0011011000;
    16'b1100000000000000: out_v[275] = 10'b1010000011;
    16'b0100000000000001: out_v[275] = 10'b0001010101;
    16'b1100000010000011: out_v[275] = 10'b0011001001;
    16'b0100000000000011: out_v[275] = 10'b1001010011;
    16'b0100000010000010: out_v[275] = 10'b1111001001;
    16'b1100000000100011: out_v[275] = 10'b0001110101;
    16'b0000000000000011: out_v[275] = 10'b1110100111;
    16'b1100010000010001: out_v[275] = 10'b0010001111;
    16'b0100010010000001: out_v[275] = 10'b0110110011;
    16'b1100010000010011: out_v[275] = 10'b1110110111;
    16'b1100010000000001: out_v[275] = 10'b1010111010;
    16'b1100000000100010: out_v[275] = 10'b1010100001;
    16'b0000100000001011: out_v[275] = 10'b0011001011;
    16'b1100000010100011: out_v[275] = 10'b1111101000;
    16'b1100000000010011: out_v[275] = 10'b1001001111;
    16'b1000000000000010: out_v[275] = 10'b1001110101;
    16'b1000000000000001: out_v[275] = 10'b0011001010;
    16'b0100000010100010: out_v[275] = 10'b1111000011;
    16'b1100000010000001: out_v[275] = 10'b1001111110;
    16'b0000000010000001: out_v[275] = 10'b0001111101;
    16'b1100010000000011: out_v[275] = 10'b0001001100;
    16'b0000010000100001: out_v[275] = 10'b1111001010;
    16'b0000000000100000: out_v[275] = 10'b0100111110;
    16'b0000000000000010: out_v[275] = 10'b1001101011;
    16'b0000000000100010: out_v[275] = 10'b1110101100;
    16'b0000000000100001: out_v[275] = 10'b0101010100;
    16'b0000000010100000: out_v[275] = 10'b1000111101;
    16'b0000000010100010: out_v[275] = 10'b0100010011;
    16'b0000000010100001: out_v[275] = 10'b1110010100;
    16'b0000000000110001: out_v[275] = 10'b1000101110;
    16'b0000000010000010: out_v[275] = 10'b1011000101;
    16'b0000000000000000: out_v[275] = 10'b0011110110;
    16'b0000010000110001: out_v[275] = 10'b1010101100;
    16'b0000010000100000: out_v[275] = 10'b1101011001;
    16'b0000000010100011: out_v[275] = 10'b0110110100;
    16'b1000000000100011: out_v[275] = 10'b1001100101;
    16'b0100000010100011: out_v[275] = 10'b0111110000;
    16'b0000000010000011: out_v[275] = 10'b0100011101;
    16'b1100000010100001: out_v[275] = 10'b0010111111;
    16'b1100010010100011: out_v[275] = 10'b1001101010;
    16'b1100000000100001: out_v[275] = 10'b1001000011;
    16'b1100100110101011: out_v[275] = 10'b0011111110;
    16'b1100100000101011: out_v[275] = 10'b1111111000;
    16'b0000100010101011: out_v[275] = 10'b0111010110;
    16'b1100000000100000: out_v[275] = 10'b0101010101;
    16'b1100100010101011: out_v[275] = 10'b1010100110;
    16'b1100000010100000: out_v[275] = 10'b0110010111;
    16'b0000010010100011: out_v[275] = 10'b1111010000;
    16'b0100000000100011: out_v[275] = 10'b1001011111;
    16'b0100100010101011: out_v[275] = 10'b1011011101;
    16'b1100000010100010: out_v[275] = 10'b0111000000;
    16'b0100010010100011: out_v[275] = 10'b1110110001;
    16'b0000100000101011: out_v[275] = 10'b0100111101;
    16'b1100100010101010: out_v[275] = 10'b0001001011;
    16'b0100000010100001: out_v[275] = 10'b0110001011;
    16'b0000000000100011: out_v[275] = 10'b1010100101;
    16'b1000000010100011: out_v[275] = 10'b0100110010;
    16'b0000100000101010: out_v[275] = 10'b0111110101;
    16'b1000000000100010: out_v[275] = 10'b1101101111;
    16'b1100100010001011: out_v[275] = 10'b0100110111;
    16'b1100000010000010: out_v[275] = 10'b0100001100;
    16'b1000000010000010: out_v[275] = 10'b0101101100;
    16'b1100000010000000: out_v[275] = 10'b1100101111;
    16'b1000000010000011: out_v[275] = 10'b0111111001;
    16'b0100000010000000: out_v[275] = 10'b0110000010;
    16'b0100010010000011: out_v[275] = 10'b0000111001;
    16'b0100000000100010: out_v[275] = 10'b0000101010;
    16'b1000000010000110: out_v[275] = 10'b1100000011;
    16'b0100000010100000: out_v[275] = 10'b1101010010;
    16'b0000000010010010: out_v[275] = 10'b0111001111;
    16'b0000000010010000: out_v[275] = 10'b1010111000;
    16'b0000000010000000: out_v[275] = 10'b0011010101;
    16'b0000010010100000: out_v[275] = 10'b1001011000;
    16'b0000000010110000: out_v[275] = 10'b1100010001;
    16'b1100000110100000: out_v[275] = 10'b0011001111;
    16'b0000010010000000: out_v[275] = 10'b1010011101;
    16'b0100010010100000: out_v[275] = 10'b0110101111;
    16'b1100010010100000: out_v[275] = 10'b1111110010;
    16'b0000000010110010: out_v[275] = 10'b0011011111;
    16'b0100000010110000: out_v[275] = 10'b0110011111;
    16'b0100000010110010: out_v[275] = 10'b1010000110;
    16'b0000000000000001: out_v[275] = 10'b1100010000;
    16'b1100000010010011: out_v[275] = 10'b1010101011;
    16'b0000000000110000: out_v[275] = 10'b0110100100;
    16'b0100000010010010: out_v[275] = 10'b0011010111;
    16'b1100010010010011: out_v[275] = 10'b1110111110;
    16'b0000000000010001: out_v[275] = 10'b0010111110;
    16'b1100000010010010: out_v[275] = 10'b0101100101;
    16'b0100000010010011: out_v[275] = 10'b0100001111;
    16'b0000000000110010: out_v[275] = 10'b1010110010;
    16'b0000000010010001: out_v[275] = 10'b1010100010;
    16'b0000000000010000: out_v[275] = 10'b0011110110;
    16'b0100000010010000: out_v[275] = 10'b0101111111;
    16'b0100010010010011: out_v[275] = 10'b0101100010;
    16'b1100010010000011: out_v[275] = 10'b0010110010;
    16'b1100010010000001: out_v[275] = 10'b1101000110;
    16'b0100000000100000: out_v[275] = 10'b0011101101;
    16'b1100010010100001: out_v[275] = 10'b1100011010;
    16'b1000000010100010: out_v[275] = 10'b1100100110;
    16'b0100010010100001: out_v[275] = 10'b1111001011;
    16'b1000000010100000: out_v[275] = 10'b1101010010;
    16'b1000000000100000: out_v[275] = 10'b1011010011;
    16'b0000000010000100: out_v[275] = 10'b0111001010;
    16'b0100000000000000: out_v[275] = 10'b0011000010;
    16'b0100000010000100: out_v[275] = 10'b1000110100;
    16'b1100000000000100: out_v[275] = 10'b1111000011;
    16'b1100000010000100: out_v[275] = 10'b0011110011;
    16'b0100000010110011: out_v[275] = 10'b0111000011;
    16'b0000000010110011: out_v[275] = 10'b1101010111;
    16'b0000000000110011: out_v[275] = 10'b1000100111;
    16'b0000000010110001: out_v[275] = 10'b0011010111;
    16'b1100000110100010: out_v[275] = 10'b1101000010;
    default: out_v[275] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1000000000000110: out_v[276] = 10'b1000110101;
    16'b1000000010100110: out_v[276] = 10'b0101010101;
    16'b0000000010100111: out_v[276] = 10'b1101000111;
    16'b1000000010100111: out_v[276] = 10'b1110010110;
    16'b1000000010000111: out_v[276] = 10'b0110011100;
    16'b0000000010100110: out_v[276] = 10'b0101001101;
    16'b0000000000100110: out_v[276] = 10'b1100110101;
    16'b1100001010100011: out_v[276] = 10'b0110100110;
    16'b1000000010000110: out_v[276] = 10'b0001010001;
    16'b1000010010100110: out_v[276] = 10'b0010001011;
    16'b1000000010100100: out_v[276] = 10'b0001011111;
    16'b1000000010100010: out_v[276] = 10'b0110000001;
    16'b0000000010000110: out_v[276] = 10'b0010100101;
    16'b1000001010100010: out_v[276] = 10'b1110100111;
    16'b1000000000100111: out_v[276] = 10'b0001001010;
    16'b1100000010100111: out_v[276] = 10'b0000110111;
    16'b1000000000100110: out_v[276] = 10'b1100110010;
    16'b1100001010100111: out_v[276] = 10'b1100011111;
    16'b0000001000100011: out_v[276] = 10'b1011100011;
    16'b0000000010100100: out_v[276] = 10'b0011010000;
    16'b0000000010100010: out_v[276] = 10'b0001000011;
    16'b1000001010100111: out_v[276] = 10'b1111000101;
    16'b1000000010100011: out_v[276] = 10'b0100000011;
    16'b0000010010100110: out_v[276] = 10'b1011000111;
    16'b1000010010000110: out_v[276] = 10'b0001011000;
    16'b1000001010100011: out_v[276] = 10'b0101110010;
    16'b1000000000100011: out_v[276] = 10'b1011011011;
    16'b1100001000100011: out_v[276] = 10'b1011100001;
    16'b1000001000100011: out_v[276] = 10'b0010011010;
    16'b1000010000000110: out_v[276] = 10'b1101000111;
    16'b1000001010100110: out_v[276] = 10'b1011011000;
    16'b0000010000000010: out_v[276] = 10'b0111000001;
    16'b0000000000000000: out_v[276] = 10'b1011010000;
    16'b0000010000000000: out_v[276] = 10'b1010001011;
    16'b1000000000000000: out_v[276] = 10'b1101000110;
    16'b1000010000000000: out_v[276] = 10'b1101101001;
    16'b1000010000000010: out_v[276] = 10'b0110000011;
    16'b0000010000100010: out_v[276] = 10'b0110100110;
    16'b0000010000100000: out_v[276] = 10'b1110100000;
    16'b1000000000000010: out_v[276] = 10'b1000110110;
    16'b0100000000000000: out_v[276] = 10'b0011010010;
    16'b1100010000000011: out_v[276] = 10'b1010110101;
    16'b1100010000000010: out_v[276] = 10'b1110111100;
    16'b1100011000000011: out_v[276] = 10'b0100000111;
    16'b1000010000100010: out_v[276] = 10'b0100110100;
    16'b1100010000100011: out_v[276] = 10'b1000000101;
    16'b0000010010100100: out_v[276] = 10'b1010011101;
    16'b1000010000100110: out_v[276] = 10'b1100111110;
    16'b1100010000100111: out_v[276] = 10'b1011011100;
    16'b1000010000100000: out_v[276] = 10'b1100110100;
    16'b1000010010100111: out_v[276] = 10'b1011001011;
    16'b1000010000100011: out_v[276] = 10'b1000000101;
    16'b1100010010100110: out_v[276] = 10'b1110101111;
    16'b1000010010100100: out_v[276] = 10'b1111010010;
    16'b1100010010100111: out_v[276] = 10'b1110110111;
    16'b1100011000100011: out_v[276] = 10'b0111011000;
    16'b1000010000000011: out_v[276] = 10'b0111110100;
    16'b1000011010100110: out_v[276] = 10'b1001101010;
    16'b1000010010100010: out_v[276] = 10'b1101110100;
    16'b1000011010100100: out_v[276] = 10'b0011101000;
    16'b1100010000000111: out_v[276] = 10'b1100110011;
    16'b1000011000100111: out_v[276] = 10'b1011011111;
    16'b1000010000100111: out_v[276] = 10'b1111011010;
    16'b1000011010100111: out_v[276] = 10'b0110100100;
    16'b1100010000100110: out_v[276] = 10'b1111000111;
    16'b0000010010100000: out_v[276] = 10'b1100010101;
    16'b1100011010100111: out_v[276] = 10'b0110101111;
    16'b1100011000100111: out_v[276] = 10'b1011101011;
    16'b1100010000100010: out_v[276] = 10'b1101110111;
    16'b0000011000000101: out_v[276] = 10'b1000010101;
    16'b1000010010100000: out_v[276] = 10'b1010010111;
    16'b1000011000100110: out_v[276] = 10'b0111111000;
    16'b1000000000000101: out_v[276] = 10'b1000011100;
    16'b1100000000000100: out_v[276] = 10'b1011011011;
    16'b1100000000000110: out_v[276] = 10'b1000011110;
    16'b1100000000000111: out_v[276] = 10'b0010111010;
    16'b0000010000000001: out_v[276] = 10'b0110011001;
    16'b1000000000000100: out_v[276] = 10'b1111100111;
    16'b1100000000100111: out_v[276] = 10'b1011110000;
    16'b0000000000000101: out_v[276] = 10'b1111011100;
    16'b1100000010000111: out_v[276] = 10'b1110111110;
    16'b1100000000000001: out_v[276] = 10'b0111001010;
    16'b1000000000000011: out_v[276] = 10'b1001000011;
    16'b1100000000100110: out_v[276] = 10'b1111111011;
    16'b1000000000100010: out_v[276] = 10'b1010111000;
    16'b1100000000000101: out_v[276] = 10'b1101110001;
    16'b1000000000000111: out_v[276] = 10'b1011011001;
    16'b0000000000000001: out_v[276] = 10'b1010000001;
    16'b1000000000000001: out_v[276] = 10'b0111101101;
    16'b0100000000000101: out_v[276] = 10'b1101100111;
    16'b1000000000100101: out_v[276] = 10'b1001001101;
    16'b0000000000000111: out_v[276] = 10'b1000111000;
    16'b1100000010000101: out_v[276] = 10'b1110100011;
    16'b0000010000000101: out_v[276] = 10'b0111100010;
    16'b1100000000000011: out_v[276] = 10'b1000011001;
    16'b0010000000000101: out_v[276] = 10'b1011010110;
    16'b1100000000000010: out_v[276] = 10'b1101010010;
    16'b1000010000000101: out_v[276] = 10'b0010101011;
    16'b0100000000000111: out_v[276] = 10'b0100001101;
    16'b1000000010000101: out_v[276] = 10'b0100001111;
    16'b0000010010000001: out_v[276] = 10'b1001110111;
    16'b0000010010000000: out_v[276] = 10'b1000100101;
    16'b0000010010000101: out_v[276] = 10'b1010010100;
    16'b0000000010000000: out_v[276] = 10'b0111110010;
    16'b0000000010000101: out_v[276] = 10'b1111100110;
    16'b1000000010000000: out_v[276] = 10'b0111100011;
    16'b0000000010000010: out_v[276] = 10'b0001101000;
    16'b0000010010000010: out_v[276] = 10'b0110011000;
    16'b0000010010000110: out_v[276] = 10'b1011111010;
    16'b0000000010000001: out_v[276] = 10'b0111000100;
    16'b0000010010000100: out_v[276] = 10'b1100011011;
    16'b0100010010000101: out_v[276] = 10'b0011110111;
    16'b0100000010000101: out_v[276] = 10'b0001011110;
    16'b1000010010000100: out_v[276] = 10'b0100110000;
    16'b0100010010100101: out_v[276] = 10'b1010110010;
    16'b0000000010000100: out_v[276] = 10'b1111000110;
    16'b0000010010100101: out_v[276] = 10'b0010110010;
    16'b1000010010000000: out_v[276] = 10'b0010111100;
    16'b1000000010000100: out_v[276] = 10'b0110011100;
    16'b0000010000000100: out_v[276] = 10'b0011001011;
    16'b0000000000000110: out_v[276] = 10'b0011101010;
    16'b0000000000100010: out_v[276] = 10'b0001011000;
    16'b0000010010100010: out_v[276] = 10'b1010011011;
    16'b0000000000000010: out_v[276] = 10'b1011001001;
    16'b0000000000000100: out_v[276] = 10'b0011100000;
    16'b0000000000100000: out_v[276] = 10'b0111100111;
    16'b1000010000000100: out_v[276] = 10'b0111011010;
    16'b0100011010000101: out_v[276] = 10'b0011101010;
    16'b0100011010000001: out_v[276] = 10'b1111000001;
    16'b1000010010000101: out_v[276] = 10'b1101111000;
    16'b0100010010100111: out_v[276] = 10'b1011100111;
    16'b0000010000000110: out_v[276] = 10'b0001101110;
    16'b1000010010000010: out_v[276] = 10'b0110111101;
    16'b0100010010000111: out_v[276] = 10'b1011111010;
    16'b1000010010000111: out_v[276] = 10'b1011101111;
    16'b0010010000000010: out_v[276] = 10'b0011010111;
    16'b0010010000000011: out_v[276] = 10'b1101000111;
    16'b0010000000000011: out_v[276] = 10'b0101101110;
    16'b0010000000000010: out_v[276] = 10'b1111110010;
    16'b0010000000000000: out_v[276] = 10'b0011100111;
    16'b0010000000000111: out_v[276] = 10'b0010100001;
    16'b0010000010000010: out_v[276] = 10'b0111101110;
    16'b0010000010000000: out_v[276] = 10'b0111010111;
    16'b0000010000000011: out_v[276] = 10'b1100110111;
    16'b0010000000000100: out_v[276] = 10'b0111011100;
    16'b0010000000000001: out_v[276] = 10'b1101110111;
    16'b0000000000000011: out_v[276] = 10'b1111011010;
    16'b1000010000100001: out_v[276] = 10'b1101101101;
    16'b1100010000000101: out_v[276] = 10'b1110010001;
    16'b1000010000000111: out_v[276] = 10'b0110000001;
    16'b1000000000100000: out_v[276] = 10'b0111110110;
    16'b1000010000000001: out_v[276] = 10'b1111010101;
    16'b0000010000000111: out_v[276] = 10'b0110101011;
    16'b0010010010000010: out_v[276] = 10'b1011001111;
    16'b0010010010000000: out_v[276] = 10'b1000100111;
    default: out_v[276] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100000000000010: out_v[277] = 10'b1011010001;
    16'b0010000001000010: out_v[277] = 10'b0000101111;
    16'b1010000001000010: out_v[277] = 10'b0111000001;
    16'b0100000001000000: out_v[277] = 10'b0001010011;
    16'b1000000001000010: out_v[277] = 10'b1001011101;
    16'b0110000001000000: out_v[277] = 10'b0101010111;
    16'b0000000000000000: out_v[277] = 10'b1100000111;
    16'b0010000000000000: out_v[277] = 10'b0100001001;
    16'b1010000001000011: out_v[277] = 10'b0101000011;
    16'b0100000001000010: out_v[277] = 10'b0010001111;
    16'b0000000001000010: out_v[277] = 10'b0101011100;
    16'b1010000000000010: out_v[277] = 10'b0010000111;
    16'b1110000001000010: out_v[277] = 10'b0010101101;
    16'b0010000001000000: out_v[277] = 10'b0001111001;
    16'b0110000001000010: out_v[277] = 10'b1011111110;
    16'b1010000001001010: out_v[277] = 10'b0100010001;
    16'b1100000001000010: out_v[277] = 10'b1000010001;
    16'b0000000001000000: out_v[277] = 10'b0101111100;
    16'b0010000000000010: out_v[277] = 10'b0011111001;
    16'b1000000001000011: out_v[277] = 10'b1111000110;
    16'b1000000000000010: out_v[277] = 10'b0110000100;
    16'b0110000101000000: out_v[277] = 10'b0100011010;
    16'b0000000000000010: out_v[277] = 10'b0010111010;
    16'b0000000100000000: out_v[277] = 10'b1000111100;
    16'b0000000101000000: out_v[277] = 10'b1010100011;
    16'b0100000101000000: out_v[277] = 10'b0001111000;
    16'b0000000101000010: out_v[277] = 10'b0101001010;
    16'b0010000100000000: out_v[277] = 10'b0111111000;
    16'b0100000100000000: out_v[277] = 10'b1101000100;
    16'b0110000100000000: out_v[277] = 10'b0000011011;
    16'b0000000100000010: out_v[277] = 10'b1100111100;
    16'b0000000101000011: out_v[277] = 10'b1010011011;
    16'b1000000101000011: out_v[277] = 10'b0010001010;
    16'b0100000101000011: out_v[277] = 10'b1011110110;
    16'b0110000100000010: out_v[277] = 10'b0100010100;
    16'b1000000101000010: out_v[277] = 10'b1011101010;
    16'b0100000100000010: out_v[277] = 10'b1100010001;
    16'b1100000101000001: out_v[277] = 10'b0101111011;
    16'b0100000101000010: out_v[277] = 10'b1101000110;
    16'b0110000101000010: out_v[277] = 10'b1010111111;
    16'b1110000101000010: out_v[277] = 10'b0101010100;
    16'b1100000101000011: out_v[277] = 10'b0100101100;
    16'b1100000100000010: out_v[277] = 10'b0001111000;
    16'b1100000100000011: out_v[277] = 10'b0011101100;
    16'b1000000100000000: out_v[277] = 10'b0100001111;
    16'b0100000001000011: out_v[277] = 10'b0110001111;
    16'b1100000100100010: out_v[277] = 10'b0001110010;
    16'b1100000101000010: out_v[277] = 10'b0010101110;
    16'b1110000100000000: out_v[277] = 10'b1110011110;
    16'b0100000101000001: out_v[277] = 10'b0001101011;
    16'b1100000101000000: out_v[277] = 10'b0110000111;
    16'b1100000001000011: out_v[277] = 10'b1000101010;
    16'b0100000101100011: out_v[277] = 10'b1011111011;
    16'b1100000101100010: out_v[277] = 10'b1010100110;
    16'b1110000100000010: out_v[277] = 10'b0110111001;
    16'b1100000100000000: out_v[277] = 10'b1100011010;
    16'b0000000001000011: out_v[277] = 10'b1010111000;
    16'b0000000100000001: out_v[277] = 10'b0011110011;
    16'b0010000101000010: out_v[277] = 10'b1001100110;
    16'b1000000100000010: out_v[277] = 10'b0001100101;
    16'b1110000101000011: out_v[277] = 10'b0010101111;
    16'b1100000100100000: out_v[277] = 10'b1001001111;
    16'b1100000101100011: out_v[277] = 10'b0111111101;
    16'b1100000000000010: out_v[277] = 10'b0010110010;
    16'b0001000101000000: out_v[277] = 10'b0101101001;
    16'b0100000000000000: out_v[277] = 10'b0111100010;
    16'b0010000101000000: out_v[277] = 10'b1101100000;
    16'b0111000101000000: out_v[277] = 10'b1110000011;
    16'b0111000100000000: out_v[277] = 10'b1101010101;
    16'b0110000000000010: out_v[277] = 10'b0011110100;
    16'b1100000100001010: out_v[277] = 10'b0101010011;
    16'b1010000101000010: out_v[277] = 10'b0001011101;
    16'b0010000100000010: out_v[277] = 10'b0001100100;
    16'b0011000101000010: out_v[277] = 10'b1000010111;
    16'b1100000000000000: out_v[277] = 10'b1111010000;
    16'b0011000001000000: out_v[277] = 10'b0011111111;
    16'b0011000101000000: out_v[277] = 10'b0100110111;
    16'b0110000000000000: out_v[277] = 10'b0000111000;
    16'b0101000101000000: out_v[277] = 10'b1100100011;
    16'b0001000100000000: out_v[277] = 10'b0011110010;
    16'b0101000001000000: out_v[277] = 10'b0111110010;
    16'b0101000100000000: out_v[277] = 10'b0010110000;
    16'b0111000001000000: out_v[277] = 10'b1111000010;
    16'b0100000000001010: out_v[277] = 10'b0011011111;
    16'b0111000101001000: out_v[277] = 10'b1011101001;
    16'b0100000001001000: out_v[277] = 10'b1110101010;
    16'b0100000100001010: out_v[277] = 10'b1000010011;
    default: out_v[277] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1000001001000011: out_v[278] = 10'b0001111100;
    16'b1100001001000011: out_v[278] = 10'b0011001101;
    16'b1100000011011011: out_v[278] = 10'b0111011111;
    16'b1000000000000011: out_v[278] = 10'b1010000011;
    16'b1100001001000010: out_v[278] = 10'b0111011011;
    16'b1100001011010010: out_v[278] = 10'b1100100101;
    16'b0100000011011001: out_v[278] = 10'b1000101110;
    16'b0000000001000011: out_v[278] = 10'b0010111001;
    16'b1100001011011010: out_v[278] = 10'b0111000100;
    16'b1100001001001010: out_v[278] = 10'b1111100100;
    16'b1100000001011011: out_v[278] = 10'b1110111110;
    16'b1100000001001001: out_v[278] = 10'b0111100101;
    16'b1100000001000011: out_v[278] = 10'b1100010111;
    16'b1000000001000001: out_v[278] = 10'b1000001111;
    16'b1100000011011001: out_v[278] = 10'b0011101101;
    16'b1100000001010001: out_v[278] = 10'b0011000011;
    16'b1100001010011010: out_v[278] = 10'b0110000001;
    16'b1000000001000011: out_v[278] = 10'b1010000111;
    16'b1100000001000010: out_v[278] = 10'b1100110111;
    16'b0100000011011110: out_v[278] = 10'b1110111100;
    16'b0100000011011101: out_v[278] = 10'b0001111110;
    16'b0100001011011001: out_v[278] = 10'b0111011111;
    16'b1100000011011010: out_v[278] = 10'b0100110000;
    16'b1100001011011011: out_v[278] = 10'b0001111111;
    16'b1100001000000010: out_v[278] = 10'b0011011101;
    16'b0100001011011110: out_v[278] = 10'b1101011011;
    16'b0100000001011001: out_v[278] = 10'b1110001100;
    16'b1100000001011001: out_v[278] = 10'b0000011111;
    16'b1100001011011001: out_v[278] = 10'b1111010111;
    16'b0100000010011101: out_v[278] = 10'b1010011111;
    16'b1100000001010011: out_v[278] = 10'b1011100100;
    16'b1100001001011011: out_v[278] = 10'b1011101111;
    16'b1100001001010011: out_v[278] = 10'b0001110111;
    16'b1100000001000001: out_v[278] = 10'b1010011011;
    16'b1100000001001011: out_v[278] = 10'b1011111010;
    16'b1100000001010010: out_v[278] = 10'b1001001110;
    16'b1100001001001001: out_v[278] = 10'b1010100111;
    16'b1000001001000010: out_v[278] = 10'b0101101110;
    16'b1100000011011101: out_v[278] = 10'b1001110111;
    16'b0100000011011100: out_v[278] = 10'b1010101110;
    16'b1100001000001010: out_v[278] = 10'b0000011011;
    16'b1100000000011001: out_v[278] = 10'b1111010100;
    16'b1100000011010011: out_v[278] = 10'b0110001010;
    16'b1000000000000001: out_v[278] = 10'b0001011010;
    16'b0100001011011101: out_v[278] = 10'b1010000101;
    16'b1100001011010011: out_v[278] = 10'b0011011011;
    16'b1010001001000011: out_v[278] = 10'b0000011011;
    16'b1100001001001011: out_v[278] = 10'b1111111110;
    16'b0010000000000000: out_v[278] = 10'b0100110011;
    16'b0010001000000000: out_v[278] = 10'b1001001100;
    16'b0000001001000001: out_v[278] = 10'b1001000011;
    16'b0010001001000000: out_v[278] = 10'b0010110001;
    16'b0010001001000001: out_v[278] = 10'b1010110111;
    16'b0000001001000000: out_v[278] = 10'b1100010001;
    16'b0000001001000011: out_v[278] = 10'b0100001000;
    16'b0010001000000001: out_v[278] = 10'b1101100000;
    16'b0000001000000010: out_v[278] = 10'b1110100110;
    16'b0000001000000000: out_v[278] = 10'b1011101101;
    16'b0010001001000011: out_v[278] = 10'b1001001011;
    16'b0000001000000001: out_v[278] = 10'b0010101010;
    16'b0000001001000010: out_v[278] = 10'b0010110011;
    16'b0000000000000000: out_v[278] = 10'b0101011111;
    16'b0010001001000010: out_v[278] = 10'b1101010100;
    16'b1100000000000010: out_v[278] = 10'b0011010110;
    16'b0000000001000010: out_v[278] = 10'b1001100011;
    16'b0010000000000001: out_v[278] = 10'b0001011100;
    16'b0010001000000010: out_v[278] = 10'b0010111111;
    16'b0010000000000010: out_v[278] = 10'b0001011101;
    16'b0110000001000010: out_v[278] = 10'b1110000110;
    16'b0010000001000001: out_v[278] = 10'b1101000100;
    16'b1000000000000010: out_v[278] = 10'b1100010110;
    16'b0110000000000010: out_v[278] = 10'b0101010100;
    16'b0000000000000010: out_v[278] = 10'b0011010110;
    16'b0010000001000000: out_v[278] = 10'b1010101100;
    16'b1010000001000010: out_v[278] = 10'b1010100010;
    16'b0010000001000010: out_v[278] = 10'b1111001001;
    16'b1110000001000010: out_v[278] = 10'b0111001000;
    16'b1110000000000010: out_v[278] = 10'b1111101000;
    16'b0110000001000000: out_v[278] = 10'b1111101110;
    16'b0110000001000110: out_v[278] = 10'b0111000110;
    16'b0010000001000011: out_v[278] = 10'b0011001010;
    16'b0110001001000010: out_v[278] = 10'b0000010100;
    16'b0000000001000000: out_v[278] = 10'b1010000011;
    16'b0100000000000010: out_v[278] = 10'b0110110010;
    16'b1000000001000010: out_v[278] = 10'b1101001100;
    16'b0110000000000000: out_v[278] = 10'b1010110101;
    16'b1110000001000000: out_v[278] = 10'b0110011101;
    16'b1010000000000010: out_v[278] = 10'b1011010011;
    16'b0000000000000001: out_v[278] = 10'b0101111010;
    16'b0000000001000001: out_v[278] = 10'b1011100110;
    16'b1110001001000010: out_v[278] = 10'b0001010100;
    16'b0010000001000110: out_v[278] = 10'b1010110111;
    16'b0010001001000110: out_v[278] = 10'b1010110111;
    16'b0110001001000110: out_v[278] = 10'b1100101101;
    16'b0000001000000011: out_v[278] = 10'b1011000010;
    16'b1000001000000010: out_v[278] = 10'b0101101011;
    16'b1000001001000001: out_v[278] = 10'b0011011010;
    16'b1010001001000001: out_v[278] = 10'b0110010000;
    16'b1000001000000011: out_v[278] = 10'b1011010111;
    16'b1000001000001001: out_v[278] = 10'b1111010011;
    16'b0000000000000011: out_v[278] = 10'b1111110001;
    16'b1000001000000001: out_v[278] = 10'b0110100000;
    16'b1000001001001001: out_v[278] = 10'b0110011010;
    16'b0010000000000011: out_v[278] = 10'b0100000010;
    16'b0010001000000011: out_v[278] = 10'b0111100010;
    16'b1010000001000011: out_v[278] = 10'b1110101000;
    16'b1010000001000001: out_v[278] = 10'b0101110011;
    16'b0110000001000011: out_v[278] = 10'b1011101110;
    16'b1010000000010010: out_v[278] = 10'b1010101111;
    16'b0110001000000000: out_v[278] = 10'b1101111000;
    16'b1110000000010010: out_v[278] = 10'b0110111010;
    16'b0000000000010010: out_v[278] = 10'b0111101110;
    16'b1110000010010010: out_v[278] = 10'b0010111011;
    16'b1010000000000000: out_v[278] = 10'b1001011101;
    16'b0110000010010011: out_v[278] = 10'b0001011111;
    16'b0110000000000011: out_v[278] = 10'b0111110010;
    16'b0110000000000001: out_v[278] = 10'b0111101001;
    16'b0110000010010010: out_v[278] = 10'b1000110001;
    16'b0010000000010010: out_v[278] = 10'b0110111011;
    16'b1110000000010000: out_v[278] = 10'b0101010011;
    16'b1110000000000000: out_v[278] = 10'b1000110110;
    16'b0110000000010010: out_v[278] = 10'b0001111011;
    16'b1110000010011000: out_v[278] = 10'b0000011010;
    16'b1110000010011010: out_v[278] = 10'b1010111001;
    16'b1110000010011011: out_v[278] = 10'b0110110111;
    16'b0010000000010011: out_v[278] = 10'b0100011011;
    16'b1110001000000000: out_v[278] = 10'b1011011001;
    16'b1110000000010011: out_v[278] = 10'b1010101011;
    16'b1110000010010000: out_v[278] = 10'b0110011011;
    16'b1010000000000011: out_v[278] = 10'b0100110110;
    16'b0110000000010011: out_v[278] = 10'b1001101111;
    16'b1110000000000001: out_v[278] = 10'b1111100110;
    16'b1010000000010011: out_v[278] = 10'b0011111010;
    16'b1110000000000011: out_v[278] = 10'b1001000110;
    16'b1110000010010011: out_v[278] = 10'b0011110101;
    16'b1100000010010010: out_v[278] = 10'b0101110111;
    16'b1010000000000001: out_v[278] = 10'b0100111011;
    16'b1000000001010001: out_v[278] = 10'b1001100111;
    16'b0000001001010011: out_v[278] = 10'b1001011011;
    16'b0010000001010011: out_v[278] = 10'b0101011010;
    16'b0100001000000000: out_v[278] = 10'b0000101101;
    16'b0000000001010001: out_v[278] = 10'b1011101010;
    16'b0000000001010011: out_v[278] = 10'b1111101110;
    16'b0100001000000010: out_v[278] = 10'b1111001010;
    16'b1000000001011001: out_v[278] = 10'b0101110111;
    16'b0010001001010011: out_v[278] = 10'b0100100110;
    16'b1000001001010001: out_v[278] = 10'b0001110010;
    16'b1010001001000010: out_v[278] = 10'b1101100011;
    16'b1110000010011110: out_v[278] = 10'b0010101011;
    16'b1110000001001010: out_v[278] = 10'b0010001111;
    16'b1010000001001010: out_v[278] = 10'b1000111110;
    16'b1110000000011010: out_v[278] = 10'b0110100110;
    16'b1000000000000000: out_v[278] = 10'b1101011001;
    16'b1100000000011010: out_v[278] = 10'b1110010010;
    16'b1110001001001010: out_v[278] = 10'b1110101011;
    16'b1110000000011110: out_v[278] = 10'b1101101011;
    16'b1010001000000010: out_v[278] = 10'b0001100010;
    16'b1010000000001010: out_v[278] = 10'b1100000111;
    16'b1010000001000000: out_v[278] = 10'b0111000011;
    16'b1010000000001000: out_v[278] = 10'b1011000111;
    16'b1000000000001000: out_v[278] = 10'b0100111001;
    16'b1100000001001010: out_v[278] = 10'b1101000111;
    16'b1010001001000000: out_v[278] = 10'b1000010110;
    16'b1110001000000010: out_v[278] = 10'b1001011111;
    16'b1110000001011010: out_v[278] = 10'b1011111000;
    16'b1000000000001010: out_v[278] = 10'b1011010110;
    16'b1100001010010011: out_v[278] = 10'b0011101110;
    16'b1000001000010010: out_v[278] = 10'b0111101010;
    16'b1000001000010011: out_v[278] = 10'b0001110000;
    16'b0001001000000010: out_v[278] = 10'b1101011001;
    16'b0000001000010000: out_v[278] = 10'b0111001101;
    16'b0000001000010001: out_v[278] = 10'b0010100011;
    16'b1000001010010011: out_v[278] = 10'b1111001010;
    16'b0000000001010000: out_v[278] = 10'b0011110111;
    16'b0000001000010011: out_v[278] = 10'b0000111111;
    16'b1000001000000000: out_v[278] = 10'b0011110011;
    16'b0001001000010010: out_v[278] = 10'b1001111011;
    16'b1001001000010010: out_v[278] = 10'b0101111111;
    16'b1000000001000000: out_v[278] = 10'b0011010110;
    16'b1000001001010011: out_v[278] = 10'b0111100010;
    16'b1010000001010011: out_v[278] = 10'b1001001111;
    16'b0010000001010001: out_v[278] = 10'b1100000011;
    16'b1010000001010001: out_v[278] = 10'b1110010110;
    16'b1110000011010010: out_v[278] = 10'b0000111111;
    16'b0110000001010011: out_v[278] = 10'b1110011011;
    16'b0110000011010011: out_v[278] = 10'b1001100111;
    16'b1110000001010011: out_v[278] = 10'b1001100101;
    16'b1100000011010010: out_v[278] = 10'b1111100110;
    16'b0110000011010010: out_v[278] = 10'b1100100111;
    16'b1010000001010010: out_v[278] = 10'b1111000110;
    16'b1110000001010010: out_v[278] = 10'b1101101111;
    16'b1000000001010011: out_v[278] = 10'b1011100110;
    16'b1110000011010011: out_v[278] = 10'b1001100011;
    16'b0001000001010010: out_v[278] = 10'b1111111111;
    16'b0000000001010010: out_v[278] = 10'b0101110101;
    16'b0011000001010010: out_v[278] = 10'b1100111111;
    16'b0010000001010010: out_v[278] = 10'b0101000111;
    16'b0011000001000010: out_v[278] = 10'b1001101011;
    16'b0110000001010010: out_v[278] = 10'b1011010011;
    16'b1110000011010000: out_v[278] = 10'b0011011111;
    16'b0010001001010010: out_v[278] = 10'b1110010001;
    default: out_v[278] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010001000000000: out_v[279] = 10'b1110001100;
    16'b0010001001111110: out_v[279] = 10'b0110001111;
    16'b0010001001001110: out_v[279] = 10'b1111000110;
    16'b1010001001001010: out_v[279] = 10'b1011110110;
    16'b0010000000000000: out_v[279] = 10'b0101100011;
    16'b0010001001001000: out_v[279] = 10'b0011001000;
    16'b0000001001001000: out_v[279] = 10'b1100001001;
    16'b0000000001001010: out_v[279] = 10'b0010010110;
    16'b0000000001001000: out_v[279] = 10'b0101001101;
    16'b0010001001001010: out_v[279] = 10'b1111010010;
    16'b0010000001001000: out_v[279] = 10'b0001011011;
    16'b0010000001001010: out_v[279] = 10'b0000011101;
    16'b1010001001001000: out_v[279] = 10'b1000101011;
    16'b0000001001001010: out_v[279] = 10'b0110001101;
    16'b0010001001011110: out_v[279] = 10'b1100101011;
    16'b0010001001011010: out_v[279] = 10'b1111101010;
    16'b0010001001101010: out_v[279] = 10'b0011100111;
    16'b1000001001001000: out_v[279] = 10'b1001100111;
    16'b0000001000000000: out_v[279] = 10'b0111001111;
    16'b0000000000000000: out_v[279] = 10'b0101110101;
    16'b1000000001001000: out_v[279] = 10'b0001100111;
    16'b0000001001101010: out_v[279] = 10'b0111001101;
    16'b0000000000100000: out_v[279] = 10'b0001101011;
    16'b0000000000010000: out_v[279] = 10'b1110100111;
    16'b0000000000110000: out_v[279] = 10'b0000111111;
    16'b0010000000000010: out_v[279] = 10'b1001111000;
    16'b0000000000000010: out_v[279] = 10'b1001011000;
    16'b0000000001011010: out_v[279] = 10'b0001011110;
    16'b0000001001011010: out_v[279] = 10'b0011111111;
    16'b0000000001011110: out_v[279] = 10'b1110011111;
    16'b0000000000001000: out_v[279] = 10'b1011101100;
    16'b1010000001001000: out_v[279] = 10'b1010110100;
    16'b0000001000100000: out_v[279] = 10'b1000101111;
    16'b0010000000100000: out_v[279] = 10'b1010100010;
    16'b0010001000000010: out_v[279] = 10'b0001011101;
    16'b0010001000100000: out_v[279] = 10'b0011011010;
    16'b0010001000100010: out_v[279] = 10'b0011001110;
    16'b0000001000000010: out_v[279] = 10'b0000111011;
    16'b0010000000100010: out_v[279] = 10'b0111000001;
    16'b0000000000100010: out_v[279] = 10'b1000111011;
    16'b0000000000000100: out_v[279] = 10'b0101111001;
    16'b0010000000010000: out_v[279] = 10'b0110101001;
    16'b0000000000010100: out_v[279] = 10'b1111100101;
    16'b0000001000000100: out_v[279] = 10'b0110001011;
    16'b0010000000010100: out_v[279] = 10'b1010100110;
    16'b0010000001011000: out_v[279] = 10'b1111010000;
    16'b0010001000000100: out_v[279] = 10'b0100110010;
    16'b0010000000000100: out_v[279] = 10'b0001011010;
    16'b1010000000000000: out_v[279] = 10'b1000010100;
    16'b0000001000010100: out_v[279] = 10'b1011101110;
    16'b0010000000001000: out_v[279] = 10'b0111010110;
    16'b0010000001011100: out_v[279] = 10'b1100011000;
    16'b0010001001001100: out_v[279] = 10'b1010100000;
    16'b0000001001001100: out_v[279] = 10'b0010101010;
    16'b0000001000000110: out_v[279] = 10'b1111000100;
    16'b0000001000010110: out_v[279] = 10'b1100100110;
    16'b0000001000110100: out_v[279] = 10'b1110001111;
    16'b0010001000010110: out_v[279] = 10'b0111000101;
    16'b0000001001011100: out_v[279] = 10'b1010110100;
    16'b0000001000010000: out_v[279] = 10'b0110111110;
    16'b0000001000100100: out_v[279] = 10'b1001110011;
    16'b0010001000010100: out_v[279] = 10'b1111010111;
    16'b0010000000010110: out_v[279] = 10'b1011001111;
    16'b0010001001011100: out_v[279] = 10'b0011010011;
    16'b0010001000000110: out_v[279] = 10'b1101101010;
    16'b0010001000001000: out_v[279] = 10'b0011100111;
    16'b0010001001011000: out_v[279] = 10'b0111011011;
    16'b1010001000000000: out_v[279] = 10'b1111011010;
    16'b0000001001101110: out_v[279] = 10'b0110100011;
    16'b0000001001011110: out_v[279] = 10'b0110100101;
    16'b0000001001111110: out_v[279] = 10'b1001011101;
    default: out_v[279] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1000000000000001: out_v[280] = 10'b1000001111;
    16'b0001001000000001: out_v[280] = 10'b1101011011;
    16'b0000000010000001: out_v[280] = 10'b1011010111;
    16'b0000000000000001: out_v[280] = 10'b0001111101;
    16'b1001000000000001: out_v[280] = 10'b1100101011;
    16'b0000000000000000: out_v[280] = 10'b0110111110;
    16'b0000100000000001: out_v[280] = 10'b0110000101;
    16'b0001000000000001: out_v[280] = 10'b1101011000;
    16'b0001100000000001: out_v[280] = 10'b1001100101;
    16'b0000001000000001: out_v[280] = 10'b0110010101;
    16'b0000001000000000: out_v[280] = 10'b0011100010;
    16'b1000001000000001: out_v[280] = 10'b1111010111;
    16'b1000000010000001: out_v[280] = 10'b1111100101;
    16'b0001000000000000: out_v[280] = 10'b1110000110;
    16'b0001001010000001: out_v[280] = 10'b1000111101;
    16'b0000001010000001: out_v[280] = 10'b1101010111;
    16'b0010010000000001: out_v[280] = 10'b0110100111;
    16'b0001000010000001: out_v[280] = 10'b0001100111;
    16'b0000100010000001: out_v[280] = 10'b1011010011;
    16'b1001001000000001: out_v[280] = 10'b0110110010;
    16'b0000000010000000: out_v[280] = 10'b1000110001;
    16'b0001001000000000: out_v[280] = 10'b0000011110;
    16'b1001000010000001: out_v[280] = 10'b0100111101;
    16'b0001010010000001: out_v[280] = 10'b0000010011;
    16'b1010010010000001: out_v[280] = 10'b0000011010;
    16'b1010010000000001: out_v[280] = 10'b1111000110;
    16'b1000000000000000: out_v[280] = 10'b1010010010;
    16'b1000010010000001: out_v[280] = 10'b0001010110;
    16'b0001000010000000: out_v[280] = 10'b1011001101;
    16'b1001000000000000: out_v[280] = 10'b1010010010;
    16'b1000010000000001: out_v[280] = 10'b1011001111;
    16'b0011010000000001: out_v[280] = 10'b1000001111;
    16'b0011010010000001: out_v[280] = 10'b0000110110;
    16'b1010000000000001: out_v[280] = 10'b1011001101;
    16'b0000010000000001: out_v[280] = 10'b1110010101;
    16'b0010000000000001: out_v[280] = 10'b1000000111;
    16'b1010000010000001: out_v[280] = 10'b0111010010;
    16'b0000010010000001: out_v[280] = 10'b1111011101;
    16'b1000000010000000: out_v[280] = 10'b1100010110;
    16'b0010010010000001: out_v[280] = 10'b0101000111;
    16'b1001001000000000: out_v[280] = 10'b0001111000;
    16'b1000001000000000: out_v[280] = 10'b1010001010;
    16'b1001001010000001: out_v[280] = 10'b1010111000;
    16'b0001001010000000: out_v[280] = 10'b1100011010;
    16'b1001000010000000: out_v[280] = 10'b1100011100;
    16'b1011010000000001: out_v[280] = 10'b0001011000;
    16'b1001000000010001: out_v[280] = 10'b0111000111;
    16'b1001001010000000: out_v[280] = 10'b0111110011;
    16'b1001010000000001: out_v[280] = 10'b1101111001;
    16'b0001100000000000: out_v[280] = 10'b1010100111;
    16'b1000000010100000: out_v[280] = 10'b0101101111;
    16'b1000010000000000: out_v[280] = 10'b1111101011;
    16'b1011000000000001: out_v[280] = 10'b1011101100;
    16'b0010000000000000: out_v[280] = 10'b0000111101;
    16'b0000010000000000: out_v[280] = 10'b0101010000;
    16'b1010010000000000: out_v[280] = 10'b0011101111;
    16'b0010010000000000: out_v[280] = 10'b0011011101;
    16'b0011000000000001: out_v[280] = 10'b1110111000;
    16'b0011000000000000: out_v[280] = 10'b1111000111;
    16'b1010000000000000: out_v[280] = 10'b1100110011;
    16'b1000010010000000: out_v[280] = 10'b1111111011;
    16'b1010010010000000: out_v[280] = 10'b1011011100;
    16'b0010010010000000: out_v[280] = 10'b1011101010;
    16'b1011010000000000: out_v[280] = 10'b1101000100;
    16'b1000000000100000: out_v[280] = 10'b0101101010;
    16'b1000100000000001: out_v[280] = 10'b1100000011;
    16'b1001100000000001: out_v[280] = 10'b1110000010;
    16'b1000101000000000: out_v[280] = 10'b0000110111;
    16'b1001101000000001: out_v[280] = 10'b0111001100;
    16'b1000101000000001: out_v[280] = 10'b0101011010;
    default: out_v[280] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000010100000: out_v[281] = 10'b0011100110;
    16'b0000010000100000: out_v[281] = 10'b1110000011;
    16'b0000010010000000: out_v[281] = 10'b0111110000;
    16'b0000110010100000: out_v[281] = 10'b0100001001;
    16'b0000100010100000: out_v[281] = 10'b0111001000;
    16'b0000000000100000: out_v[281] = 10'b0010011110;
    16'b0000010000000000: out_v[281] = 10'b0001111011;
    16'b0000100010000000: out_v[281] = 10'b0110111011;
    16'b0000010010100000: out_v[281] = 10'b1110010001;
    16'b0000000010000000: out_v[281] = 10'b0000111011;
    16'b0000110010000000: out_v[281] = 10'b0101100010;
    16'b0000110000100000: out_v[281] = 10'b0000110101;
    16'b0000000000000000: out_v[281] = 10'b1001010101;
    16'b0000100000000000: out_v[281] = 10'b0000101110;
    16'b0000100000100000: out_v[281] = 10'b0000001100;
    16'b0000000000010000: out_v[281] = 10'b0000000110;
    16'b0000100000000010: out_v[281] = 10'b0111010110;
    16'b0001000000000000: out_v[281] = 10'b1111001011;
    16'b0000110000000000: out_v[281] = 10'b1101111010;
    16'b0000010000000100: out_v[281] = 10'b1011100100;
    16'b0000000000000100: out_v[281] = 10'b1110000000;
    16'b0000000110000000: out_v[281] = 10'b1010000011;
    16'b0000000100000000: out_v[281] = 10'b1111001000;
    16'b0000010010000100: out_v[281] = 10'b1111111000;
    16'b0000000010000100: out_v[281] = 10'b0111111010;
    default: out_v[281] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1000110000000000: out_v[282] = 10'b0001110001;
    16'b1000110001000000: out_v[282] = 10'b1011110110;
    16'b1100100001100000: out_v[282] = 10'b0110001011;
    16'b0000010000100000: out_v[282] = 10'b0101000101;
    16'b0000010000000000: out_v[282] = 10'b1100000101;
    16'b0000000000100000: out_v[282] = 10'b1010010001;
    16'b1000100001000000: out_v[282] = 10'b0010001110;
    16'b0100010001100000: out_v[282] = 10'b1000001110;
    16'b0100000001000000: out_v[282] = 10'b1001001011;
    16'b1000110001100000: out_v[282] = 10'b1010100001;
    16'b1000110000001000: out_v[282] = 10'b0111010010;
    16'b1100110001100000: out_v[282] = 10'b0111101011;
    16'b0000000000000000: out_v[282] = 10'b0110110000;
    16'b0000010001000000: out_v[282] = 10'b0101100110;
    16'b1000100000000000: out_v[282] = 10'b0010110010;
    16'b0100000001100000: out_v[282] = 10'b1101001011;
    16'b1000110000100000: out_v[282] = 10'b1011100010;
    16'b0100010000100000: out_v[282] = 10'b0010111010;
    16'b0000010001100000: out_v[282] = 10'b1000110011;
    16'b0000010000100010: out_v[282] = 10'b1000010101;
    16'b0000110000000000: out_v[282] = 10'b1001110100;
    16'b1000010000000000: out_v[282] = 10'b1101100101;
    16'b1000100001100000: out_v[282] = 10'b1111010100;
    16'b0000110000100000: out_v[282] = 10'b0101110000;
    16'b0100010001000000: out_v[282] = 10'b0010001011;
    16'b0100110001100000: out_v[282] = 10'b1100111110;
    16'b0000000001100000: out_v[282] = 10'b1001011111;
    16'b0000110001100000: out_v[282] = 10'b1110110110;
    16'b0000000000001000: out_v[282] = 10'b0011001010;
    16'b1000010000001000: out_v[282] = 10'b0010001110;
    16'b0000010000001000: out_v[282] = 10'b1000101000;
    16'b1000000000001000: out_v[282] = 10'b1000101111;
    16'b1000100000001000: out_v[282] = 10'b1001110110;
    16'b0000000000001010: out_v[282] = 10'b0011111101;
    16'b0001010000001010: out_v[282] = 10'b1010011111;
    16'b0000000000000010: out_v[282] = 10'b0001100010;
    16'b0000010000000010: out_v[282] = 10'b1010100111;
    16'b0000010000001010: out_v[282] = 10'b1001100101;
    16'b0001010000000000: out_v[282] = 10'b0011010110;
    16'b0001010000000010: out_v[282] = 10'b1100101110;
    16'b1000010000001010: out_v[282] = 10'b1000100110;
    16'b0000010000101000: out_v[282] = 10'b1010010001;
    16'b0001000000000010: out_v[282] = 10'b0000100111;
    16'b0001000000001010: out_v[282] = 10'b0011011001;
    16'b0000000001000000: out_v[282] = 10'b1110010110;
    16'b1000110000001010: out_v[282] = 10'b0100011001;
    16'b1000000000001010: out_v[282] = 10'b0011111100;
    16'b1000100000001010: out_v[282] = 10'b1100110010;
    16'b1000110000101000: out_v[282] = 10'b1001001011;
    16'b1000110000101010: out_v[282] = 10'b0111011011;
    16'b1000000000000000: out_v[282] = 10'b1101011000;
    16'b1000100000000010: out_v[282] = 10'b1010001100;
    16'b1001110000001010: out_v[282] = 10'b0000110111;
    16'b1001010000001010: out_v[282] = 10'b0000101010;
    16'b1000110000000010: out_v[282] = 10'b0110110110;
    16'b1001100000001010: out_v[282] = 10'b1011001010;
    16'b0000000000101000: out_v[282] = 10'b1011110010;
    16'b0000100000000000: out_v[282] = 10'b0110111000;
    16'b0100000000100000: out_v[282] = 10'b0100010111;
    16'b1000100000100000: out_v[282] = 10'b0001111010;
    16'b1000100001001000: out_v[282] = 10'b0000110010;
    16'b1000000001001000: out_v[282] = 10'b0110001011;
    16'b0000100001000000: out_v[282] = 10'b0100101110;
    16'b1000010000101000: out_v[282] = 10'b0100110110;
    16'b1000000001000000: out_v[282] = 10'b1000100001;
    16'b0000000000100010: out_v[282] = 10'b1111000011;
    16'b0000000000101010: out_v[282] = 10'b1110111000;
    16'b1000100000101000: out_v[282] = 10'b0110001011;
    16'b1000110001001000: out_v[282] = 10'b0111110000;
    16'b1000010001001000: out_v[282] = 10'b0110110110;
    16'b0000010001001000: out_v[282] = 10'b1100001000;
    16'b0000110000001000: out_v[282] = 10'b0111110001;
    16'b0000000001001000: out_v[282] = 10'b1100011011;
    16'b0000100000001000: out_v[282] = 10'b1101001110;
    default: out_v[282] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001011000000100: out_v[283] = 10'b1001110111;
    16'b0001100000000100: out_v[283] = 10'b0101001100;
    16'b0001010000000100: out_v[283] = 10'b0000110001;
    16'b0101010000000100: out_v[283] = 10'b0100110001;
    16'b0000010000000100: out_v[283] = 10'b1000011101;
    16'b0001000000000000: out_v[283] = 10'b0010110101;
    16'b0000010000000000: out_v[283] = 10'b0110001110;
    16'b0001000000000100: out_v[283] = 10'b0010001001;
    16'b0001010000000000: out_v[283] = 10'b0011011001;
    16'b0001000000001100: out_v[283] = 10'b0011101000;
    16'b0001110000000100: out_v[283] = 10'b1110100000;
    16'b0100010000000100: out_v[283] = 10'b0011000001;
    16'b0000000000000100: out_v[283] = 10'b1000111100;
    16'b0000011000000100: out_v[283] = 10'b1001101101;
    16'b0000000000001100: out_v[283] = 10'b0101000101;
    16'b0100011000000100: out_v[283] = 10'b0110010111;
    16'b0101010000000000: out_v[283] = 10'b0110011110;
    16'b0001001000000100: out_v[283] = 10'b0000011001;
    16'b0011010000000100: out_v[283] = 10'b0011011011;
    16'b0001011000001100: out_v[283] = 10'b1011110110;
    16'b0001010000001100: out_v[283] = 10'b0101100110;
    16'b0010000000001100: out_v[283] = 10'b0110101000;
    16'b0010001000000000: out_v[283] = 10'b1101010011;
    16'b0010000000000000: out_v[283] = 10'b1101000111;
    16'b0010000000001000: out_v[283] = 10'b0100110110;
    16'b0010000000000100: out_v[283] = 10'b1101000100;
    16'b0010100000001000: out_v[283] = 10'b1110000001;
    16'b0000000000001000: out_v[283] = 10'b1101010000;
    16'b0010001000001000: out_v[283] = 10'b0111001011;
    16'b0010100000001100: out_v[283] = 10'b1111110010;
    16'b0010001000001100: out_v[283] = 10'b1110100010;
    16'b0010000001001000: out_v[283] = 10'b1010011111;
    16'b0000000000000000: out_v[283] = 10'b1111101010;
    16'b0010010000001000: out_v[283] = 10'b0010001111;
    16'b0011000000001000: out_v[283] = 10'b0100100100;
    16'b0010010000001100: out_v[283] = 10'b0010001100;
    16'b0010010000000100: out_v[283] = 10'b0011011110;
    16'b0110000000000000: out_v[283] = 10'b1100010111;
    16'b0110000000001000: out_v[283] = 10'b0011010101;
    16'b0111000000001000: out_v[283] = 10'b1010100111;
    16'b0011000000001100: out_v[283] = 10'b1000101100;
    16'b0011000000000000: out_v[283] = 10'b1111000001;
    16'b0010010000000000: out_v[283] = 10'b1111000000;
    16'b0011010000001000: out_v[283] = 10'b1101011001;
    16'b0010001000000100: out_v[283] = 10'b1101010111;
    16'b0011010000001100: out_v[283] = 10'b1100110011;
    16'b0000001000000100: out_v[283] = 10'b1001011101;
    16'b0011001000001100: out_v[283] = 10'b1100101000;
    16'b0010001010001000: out_v[283] = 10'b0011011001;
    16'b0001100000001100: out_v[283] = 10'b1000101011;
    16'b0001001000001100: out_v[283] = 10'b0110101111;
    16'b0100000000000100: out_v[283] = 10'b0111111001;
    16'b0000001000001100: out_v[283] = 10'b1111110111;
    16'b0010011000001100: out_v[283] = 10'b0011001011;
    16'b0000100000000100: out_v[283] = 10'b0111011011;
    16'b0000100000001100: out_v[283] = 10'b0100110011;
    16'b0011100000001100: out_v[283] = 10'b1000111110;
    16'b0000001000000000: out_v[283] = 10'b1001011100;
    16'b0010110000001100: out_v[283] = 10'b0011001101;
    16'b0000010000001100: out_v[283] = 10'b0110011110;
    16'b0001001000000000: out_v[283] = 10'b1110111000;
    16'b0001010000001000: out_v[283] = 10'b1001000011;
    16'b0011011010001000: out_v[283] = 10'b1001100111;
    16'b0001011010001000: out_v[283] = 10'b1100110111;
    16'b0001000000001000: out_v[283] = 10'b1101011011;
    16'b0011011000001000: out_v[283] = 10'b1001111001;
    16'b0011001000001000: out_v[283] = 10'b0110010001;
    16'b0001011000000000: out_v[283] = 10'b1011111100;
    16'b0011010000000000: out_v[283] = 10'b1001011000;
    16'b0011000000001101: out_v[283] = 10'b1011101111;
    16'b0010011000001000: out_v[283] = 10'b0110111000;
    16'b0011011000000000: out_v[283] = 10'b1010111100;
    16'b0011000000000100: out_v[283] = 10'b0011000110;
    16'b0001011000001000: out_v[283] = 10'b1001100010;
    16'b0111010000001000: out_v[283] = 10'b1011111010;
    16'b0011001010001000: out_v[283] = 10'b1001010101;
    16'b0011010000001101: out_v[283] = 10'b1010010101;
    16'b0011001000000000: out_v[283] = 10'b0111001011;
    16'b0001011000000101: out_v[283] = 10'b1010011000;
    16'b0011011000001100: out_v[283] = 10'b0100110010;
    16'b0001010001000100: out_v[283] = 10'b0100110110;
    16'b0001000000000101: out_v[283] = 10'b1101011110;
    16'b0011011000001101: out_v[283] = 10'b1011001100;
    16'b0001000000001101: out_v[283] = 10'b0111010111;
    16'b0001010000000101: out_v[283] = 10'b0100011110;
    16'b0010000000001101: out_v[283] = 10'b1011011001;
    16'b0011100000001101: out_v[283] = 10'b0101111101;
    16'b0001111000000100: out_v[283] = 10'b0110100110;
    16'b1011000000001000: out_v[283] = 10'b1110100111;
    16'b1011010000001000: out_v[283] = 10'b1111101000;
    16'b1011000000000000: out_v[283] = 10'b1101001011;
    16'b1001000000000000: out_v[283] = 10'b1011010100;
    16'b1010000000001000: out_v[283] = 10'b0111001101;
    16'b1011010000000000: out_v[283] = 10'b0101111101;
    16'b1000000000001000: out_v[283] = 10'b1111111000;
    16'b1001000000001000: out_v[283] = 10'b0110110111;
    16'b1010000000000000: out_v[283] = 10'b1010001111;
    16'b0010110000000100: out_v[283] = 10'b0011110111;
    16'b0000011010000000: out_v[283] = 10'b1111100010;
    16'b0010011010001000: out_v[283] = 10'b0011101011;
    16'b0000001010000000: out_v[283] = 10'b0010011011;
    16'b0010011010000000: out_v[283] = 10'b1111100011;
    16'b0000110000000100: out_v[283] = 10'b0111011110;
    16'b0001011010000000: out_v[283] = 10'b0111001100;
    16'b0011011010000000: out_v[283] = 10'b1011001000;
    16'b0000011000000000: out_v[283] = 10'b1001100111;
    16'b0010011000000000: out_v[283] = 10'b1101100011;
    16'b0010100000000100: out_v[283] = 10'b1001110011;
    16'b0010011000000100: out_v[283] = 10'b0110100101;
    16'b0010011010000100: out_v[283] = 10'b0101010110;
    16'b0011110000000100: out_v[283] = 10'b0010001110;
    16'b0010001010000000: out_v[283] = 10'b1110000100;
    16'b0011110000001100: out_v[283] = 10'b1001100011;
    16'b0011011010001100: out_v[283] = 10'b0111100101;
    16'b0000011000001100: out_v[283] = 10'b0111110111;
    16'b0011011000000100: out_v[283] = 10'b0100001011;
    16'b0010100000001101: out_v[283] = 10'b1110000101;
    16'b0011001010000000: out_v[283] = 10'b1001001011;
    16'b0001001010001000: out_v[283] = 10'b1111000100;
    16'b0000010000001000: out_v[283] = 10'b1111000110;
    16'b0000011010001000: out_v[283] = 10'b1001111110;
    default: out_v[283] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000011000001010: out_v[284] = 10'b1100001011;
    16'b0000111000000010: out_v[284] = 10'b0000000101;
    16'b0000110000000010: out_v[284] = 10'b0111111010;
    16'b0000101000000010: out_v[284] = 10'b1011110010;
    16'b0000110000001010: out_v[284] = 10'b1101100000;
    16'b0000001000000010: out_v[284] = 10'b1001010101;
    16'b0000110000000000: out_v[284] = 10'b0010100110;
    16'b0000100000000010: out_v[284] = 10'b1011100011;
    16'b0000011000000010: out_v[284] = 10'b0100100101;
    16'b0100111000001010: out_v[284] = 10'b0101000000;
    16'b0000111000001010: out_v[284] = 10'b0001110001;
    16'b0000101000001010: out_v[284] = 10'b0100011011;
    16'b0000010000000010: out_v[284] = 10'b0011010001;
    16'b0000010000000000: out_v[284] = 10'b0111100011;
    16'b0000101000000000: out_v[284] = 10'b1010101001;
    16'b0000010000001000: out_v[284] = 10'b0110111001;
    16'b0100011000001010: out_v[284] = 10'b0001001111;
    16'b0000010000001010: out_v[284] = 10'b1110100111;
    16'b0000110000001000: out_v[284] = 10'b0110110110;
    16'b0000101000001000: out_v[284] = 10'b0010011101;
    16'b0100011000001000: out_v[284] = 10'b1001111010;
    16'b0100010000000000: out_v[284] = 10'b0001111011;
    16'b0100000000000000: out_v[284] = 10'b1100010111;
    16'b0100000000001000: out_v[284] = 10'b1100001011;
    16'b0100010000001000: out_v[284] = 10'b0000101101;
    16'b0100011000000000: out_v[284] = 10'b1011110100;
    16'b0100011000000010: out_v[284] = 10'b0110110000;
    16'b0100100000001000: out_v[284] = 10'b1100010110;
    16'b0100100000000000: out_v[284] = 10'b1111000101;
    16'b0110000000000000: out_v[284] = 10'b1101100101;
    16'b0110011000001010: out_v[284] = 10'b1110000110;
    16'b0100010000001010: out_v[284] = 10'b1000101110;
    16'b0000001000000000: out_v[284] = 10'b1001011011;
    16'b0000011000000000: out_v[284] = 10'b1000101100;
    16'b0100001000001000: out_v[284] = 10'b0011000100;
    16'b0000000000000000: out_v[284] = 10'b1000000000;
    16'b0100001000001010: out_v[284] = 10'b1011101110;
    16'b0010001000000010: out_v[284] = 10'b1110110011;
    16'b0100001000000010: out_v[284] = 10'b0001011010;
    16'b0000001000001010: out_v[284] = 10'b0111011000;
    16'b0000000000000010: out_v[284] = 10'b1001001101;
    16'b0010011000000010: out_v[284] = 10'b0000000001;
    16'b0100101000001010: out_v[284] = 10'b0001111010;
    16'b0100111000000010: out_v[284] = 10'b0011110101;
    16'b0000100000000000: out_v[284] = 10'b0111001101;
    16'b0100101000000010: out_v[284] = 10'b1001100110;
    16'b0110011000000010: out_v[284] = 10'b0001110111;
    16'b0110001000000010: out_v[284] = 10'b1111110010;
    16'b0010111000000010: out_v[284] = 10'b0111000101;
    16'b0110001000001010: out_v[284] = 10'b0110011010;
    16'b0010010000000000: out_v[284] = 10'b1011010100;
    16'b0100110000001010: out_v[284] = 10'b0011011010;
    16'b0000000000001000: out_v[284] = 10'b0111010001;
    16'b0100000001001000: out_v[284] = 10'b1001011111;
    16'b0110010000001000: out_v[284] = 10'b1110011010;
    16'b0100100001001000: out_v[284] = 10'b1100000101;
    16'b0100110000001000: out_v[284] = 10'b1001110000;
    16'b0100010000000010: out_v[284] = 10'b0001011001;
    16'b0100110000000000: out_v[284] = 10'b0111000011;
    16'b0000100000001000: out_v[284] = 10'b0111000011;
    16'b0010000000000000: out_v[284] = 10'b0000010100;
    16'b0000000001001000: out_v[284] = 10'b0101011000;
    16'b0000000001000000: out_v[284] = 10'b0001101111;
    16'b0000001000001000: out_v[284] = 10'b0011100100;
    16'b0000100001001000: out_v[284] = 10'b0111001110;
    16'b0100101000001000: out_v[284] = 10'b1101001110;
    16'b0100101000000000: out_v[284] = 10'b0011110011;
    16'b0000100001000000: out_v[284] = 10'b0001000100;
    16'b0100000000001010: out_v[284] = 10'b0100101100;
    16'b0100100000001010: out_v[284] = 10'b1100101111;
    16'b0100111000001000: out_v[284] = 10'b0111111000;
    16'b0000000000001010: out_v[284] = 10'b0101101000;
    16'b0000011000001000: out_v[284] = 10'b0001110111;
    16'b0100001000000000: out_v[284] = 10'b0011111000;
    16'b0001100001000000: out_v[284] = 10'b0111010010;
    16'b0100100001000000: out_v[284] = 10'b0011100101;
    16'b0000101001000000: out_v[284] = 10'b1101111111;
    16'b0100000001000000: out_v[284] = 10'b1110100100;
    16'b0001100000000000: out_v[284] = 10'b1011000011;
    16'b0110000000001000: out_v[284] = 10'b0100110001;
    16'b0000111000001000: out_v[284] = 10'b0000111011;
    16'b0000101001000010: out_v[284] = 10'b1111000000;
    16'b0100101001000000: out_v[284] = 10'b0101010101;
    default: out_v[284] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1000010000000000: out_v[285] = 10'b0100110011;
    16'b1000011000000000: out_v[285] = 10'b0000011001;
    16'b1000101000000000: out_v[285] = 10'b1111001100;
    16'b1000100000000000: out_v[285] = 10'b1000100110;
    16'b1000001000000000: out_v[285] = 10'b1001001101;
    16'b0000000000000000: out_v[285] = 10'b1110000011;
    16'b1000100000010000: out_v[285] = 10'b0000110001;
    16'b1000111000010000: out_v[285] = 10'b1010110001;
    16'b0000010000000000: out_v[285] = 10'b1101100101;
    16'b0000011000000000: out_v[285] = 10'b0000111101;
    16'b0000001000000000: out_v[285] = 10'b0001110101;
    16'b1000000000000000: out_v[285] = 10'b0100000111;
    16'b1000000000010000: out_v[285] = 10'b1011001101;
    16'b1000010000010000: out_v[285] = 10'b1010001011;
    16'b1000110000010000: out_v[285] = 10'b0110100010;
    16'b1000101000010000: out_v[285] = 10'b1110110101;
    16'b0000100000010000: out_v[285] = 10'b1001110100;
    16'b0000100000000000: out_v[285] = 10'b0001001101;
    16'b1000110000000000: out_v[285] = 10'b0100110010;
    16'b1000111000000000: out_v[285] = 10'b0110001111;
    16'b1000011000010000: out_v[285] = 10'b0010110111;
    16'b1000100100010000: out_v[285] = 10'b1000110101;
    16'b0000000000010000: out_v[285] = 10'b1011011100;
    16'b0000001000010000: out_v[285] = 10'b0100011110;
    16'b1000000000010010: out_v[285] = 10'b1010011111;
    16'b0000011000010000: out_v[285] = 10'b0001101101;
    16'b1000001000010000: out_v[285] = 10'b0111001000;
    16'b1000001100010000: out_v[285] = 10'b1000011000;
    16'b1000011000100000: out_v[285] = 10'b0010011101;
    16'b0000000000010010: out_v[285] = 10'b0111011101;
    16'b1000000100010000: out_v[285] = 10'b1110001100;
    16'b1000001000010010: out_v[285] = 10'b0111000111;
    16'b1000011000010010: out_v[285] = 10'b0110111111;
    16'b1000101100010000: out_v[285] = 10'b1101000100;
    16'b0000101000000000: out_v[285] = 10'b1000011111;
    16'b0000010000010000: out_v[285] = 10'b1000111100;
    16'b1000011000000010: out_v[285] = 10'b0011100110;
    16'b1000010100010000: out_v[285] = 10'b1101001011;
    16'b1000111100010000: out_v[285] = 10'b0001001110;
    16'b1000011100010000: out_v[285] = 10'b1000010100;
    16'b0000010100010000: out_v[285] = 10'b1110011010;
    16'b0001011000000000: out_v[285] = 10'b1111010111;
    16'b0000111000000000: out_v[285] = 10'b0011100100;
    16'b0000111000010000: out_v[285] = 10'b1011100110;
    16'b0010010000000000: out_v[285] = 10'b0011111111;
    16'b0000101000010000: out_v[285] = 10'b1011000001;
    16'b0001011000000001: out_v[285] = 10'b0011111000;
    16'b1000111100000010: out_v[285] = 10'b0001110100;
    16'b1000111100000000: out_v[285] = 10'b0111010001;
    16'b1010011000000000: out_v[285] = 10'b1111001010;
    16'b1001010000000001: out_v[285] = 10'b1101100001;
    16'b1001011000000001: out_v[285] = 10'b1011100110;
    16'b0000110000010000: out_v[285] = 10'b1011110010;
    16'b1001000000000000: out_v[285] = 10'b0111111100;
    16'b1010101100000000: out_v[285] = 10'b1111011001;
    16'b1001001000000001: out_v[285] = 10'b1101101100;
    16'b0000101100000000: out_v[285] = 10'b0010000011;
    16'b1001100000000000: out_v[285] = 10'b0011111101;
    16'b0001001000000000: out_v[285] = 10'b1011100100;
    16'b1010000000000000: out_v[285] = 10'b1010111001;
    16'b1001101000000001: out_v[285] = 10'b0111110011;
    16'b0001000000000000: out_v[285] = 10'b0111001101;
    16'b0000001100000000: out_v[285] = 10'b1001100110;
    16'b1001101000000000: out_v[285] = 10'b1001011011;
    16'b0001101100000001: out_v[285] = 10'b1011011000;
    16'b1000101100000000: out_v[285] = 10'b0111000011;
    16'b0010101000000000: out_v[285] = 10'b1010011110;
    16'b1000101100000001: out_v[285] = 10'b1101110011;
    16'b1001100000000001: out_v[285] = 10'b1011111110;
    16'b0001101000000001: out_v[285] = 10'b0011111010;
    16'b1010101000000000: out_v[285] = 10'b0011101111;
    16'b1001011000000000: out_v[285] = 10'b1101100110;
    16'b1010001000000000: out_v[285] = 10'b1001110011;
    16'b1000101000000001: out_v[285] = 10'b1001111011;
    16'b1001101100000001: out_v[285] = 10'b1001111001;
    16'b0001001000000001: out_v[285] = 10'b1111001110;
    16'b1000001100000000: out_v[285] = 10'b0110010011;
    16'b0001101000000000: out_v[285] = 10'b0111011011;
    16'b1010100000000000: out_v[285] = 10'b1011110001;
    16'b0000001010000000: out_v[285] = 10'b0110101101;
    16'b0000001011000000: out_v[285] = 10'b1101101110;
    16'b1001111000000001: out_v[285] = 10'b1110000110;
    16'b1001101100000000: out_v[285] = 10'b1111110011;
    16'b0010001000000000: out_v[285] = 10'b1111100111;
    16'b0010000000000000: out_v[285] = 10'b0110110111;
    16'b1001001000000000: out_v[285] = 10'b1101111010;
    16'b1001010000000000: out_v[285] = 10'b1111000010;
    16'b0000101011000000: out_v[285] = 10'b0001111111;
    16'b1001000000000001: out_v[285] = 10'b0111010011;
    16'b0001101100000000: out_v[285] = 10'b0111110101;
    16'b1001001100000001: out_v[285] = 10'b1001111101;
    16'b1010010000000000: out_v[285] = 10'b1100000111;
    16'b0000101000000001: out_v[285] = 10'b1101110110;
    16'b0000101100000001: out_v[285] = 10'b1111011001;
    16'b0000101110000000: out_v[285] = 10'b0010110110;
    16'b1000011000000001: out_v[285] = 10'b1101100100;
    16'b1000010000000001: out_v[285] = 10'b1111010101;
    16'b1001111000000000: out_v[285] = 10'b1101100110;
    16'b1000001000000001: out_v[285] = 10'b0111000001;
    default: out_v[285] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1000100010000100: out_v[286] = 10'b1000101010;
    16'b1100110110000100: out_v[286] = 10'b1111001001;
    16'b0100100010000100: out_v[286] = 10'b0011011010;
    16'b0000100010000100: out_v[286] = 10'b0000111100;
    16'b1000100000000100: out_v[286] = 10'b0100111001;
    16'b0000100000000110: out_v[286] = 10'b0001001011;
    16'b0000100000000000: out_v[286] = 10'b1100000110;
    16'b0100000010000100: out_v[286] = 10'b0100110110;
    16'b0000000010000100: out_v[286] = 10'b0100001001;
    16'b1100000010000100: out_v[286] = 10'b0111100010;
    16'b0000000000000100: out_v[286] = 10'b1101100110;
    16'b1100100000000100: out_v[286] = 10'b0010110001;
    16'b1100010110000100: out_v[286] = 10'b0111100011;
    16'b0000100110000100: out_v[286] = 10'b0011011111;
    16'b0100000010001100: out_v[286] = 10'b1000101101;
    16'b1000000010000100: out_v[286] = 10'b0101101100;
    16'b0000100000000100: out_v[286] = 10'b0000101101;
    16'b1100100010000100: out_v[286] = 10'b0001011010;
    16'b0000100010000110: out_v[286] = 10'b0001000001;
    16'b1100100010001100: out_v[286] = 10'b0011110111;
    16'b1100100000001100: out_v[286] = 10'b0110011011;
    16'b1000100010000110: out_v[286] = 10'b0110011011;
    16'b1000100110000100: out_v[286] = 10'b0101101001;
    16'b0000100000000010: out_v[286] = 10'b0001100111;
    16'b1100100000000101: out_v[286] = 10'b0110001011;
    16'b0100110110000100: out_v[286] = 10'b1110100101;
    16'b0000100010000000: out_v[286] = 10'b1110000001;
    16'b0100100110000100: out_v[286] = 10'b1101110101;
    16'b1100000010001100: out_v[286] = 10'b0100101011;
    16'b1000100010000000: out_v[286] = 10'b0110110011;
    16'b1000100000000101: out_v[286] = 10'b0111001001;
    16'b0100100010000110: out_v[286] = 10'b1100000111;
    16'b1100100110000100: out_v[286] = 10'b0111001001;
    16'b0000000010000110: out_v[286] = 10'b1010010011;
    16'b1100110110000000: out_v[286] = 10'b1100000001;
    16'b0100100000001100: out_v[286] = 10'b0010010110;
    16'b0000100100000100: out_v[286] = 10'b1100101101;
    16'b0000000010000000: out_v[286] = 10'b1010100111;
    16'b1000000000000000: out_v[286] = 10'b0101000110;
    16'b0000000000000000: out_v[286] = 10'b0011010100;
    16'b1000000010000000: out_v[286] = 10'b0010111011;
    16'b0100100000000100: out_v[286] = 10'b0101010100;
    16'b0100110000000100: out_v[286] = 10'b0011010010;
    16'b0100110100000100: out_v[286] = 10'b1011000001;
    16'b0000100000001100: out_v[286] = 10'b1010111011;
    16'b0000000100000000: out_v[286] = 10'b0011111011;
    16'b0000100100000000: out_v[286] = 10'b1111100000;
    16'b0000100110000000: out_v[286] = 10'b1010010010;
    16'b0000000000000110: out_v[286] = 10'b0011011010;
    16'b0100100000000110: out_v[286] = 10'b1000110001;
    16'b0000000000000010: out_v[286] = 10'b1001000100;
    16'b0000000000001101: out_v[286] = 10'b0100011110;
    16'b0000100000000111: out_v[286] = 10'b0111111011;
    16'b0000100000000001: out_v[286] = 10'b1000000110;
    16'b0000100000000101: out_v[286] = 10'b1100011011;
    16'b1000000000000100: out_v[286] = 10'b1011100010;
    16'b1000100000000110: out_v[286] = 10'b0010000110;
    16'b0100000000000100: out_v[286] = 10'b0100010111;
    16'b0000000000001100: out_v[286] = 10'b1001100101;
    16'b1000000000000110: out_v[286] = 10'b1100111100;
    16'b1000000000000010: out_v[286] = 10'b0101101011;
    16'b0000100000001101: out_v[286] = 10'b0010111110;
    16'b1000100000000000: out_v[286] = 10'b0000110001;
    16'b0000000000000101: out_v[286] = 10'b0111101110;
    16'b1100010110000000: out_v[286] = 10'b1000110010;
    16'b0100110110000000: out_v[286] = 10'b0000111110;
    16'b1000100110000000: out_v[286] = 10'b1010100110;
    16'b1100100010000000: out_v[286] = 10'b1011101100;
    16'b1000000110000000: out_v[286] = 10'b1100011011;
    16'b1000000010000010: out_v[286] = 10'b0001101110;
    16'b1100100010000101: out_v[286] = 10'b0101110111;
    16'b0100100010000101: out_v[286] = 10'b1111110000;
    16'b1100100010001101: out_v[286] = 10'b1010100110;
    16'b1100000010000000: out_v[286] = 10'b1011101100;
    16'b0100010110000000: out_v[286] = 10'b0101000011;
    16'b1000000010000110: out_v[286] = 10'b1001110111;
    16'b1000100100000000: out_v[286] = 10'b1001011100;
    16'b1000100010001000: out_v[286] = 10'b1100110100;
    16'b0000000110000000: out_v[286] = 10'b1011010010;
    16'b1000000100000000: out_v[286] = 10'b0010011000;
    16'b0000100010001000: out_v[286] = 10'b0010110010;
    16'b1100010100000100: out_v[286] = 10'b0101110101;
    16'b0000000010001000: out_v[286] = 10'b0100111000;
    16'b0000000000001000: out_v[286] = 10'b0110101100;
    16'b1100010000000100: out_v[286] = 10'b0010110100;
    16'b0000100000001000: out_v[286] = 10'b1110011000;
    16'b1000100000001000: out_v[286] = 10'b1101000010;
    16'b1100000110000100: out_v[286] = 10'b0011001101;
    16'b1000000000001100: out_v[286] = 10'b0101100101;
    16'b1000000010001100: out_v[286] = 10'b1010100100;
    16'b1000100010001100: out_v[286] = 10'b1101011101;
    16'b1000000110000100: out_v[286] = 10'b1110011100;
    16'b1000100000001100: out_v[286] = 10'b1101000100;
    16'b1000000000001000: out_v[286] = 10'b0110000011;
    16'b0000110100000000: out_v[286] = 10'b0111110101;
    16'b0000100001000000: out_v[286] = 10'b0011011111;
    16'b0100110100000000: out_v[286] = 10'b0011001011;
    16'b1100110100000100: out_v[286] = 10'b1010100110;
    16'b0000110110000000: out_v[286] = 10'b0001101101;
    16'b1000110110000000: out_v[286] = 10'b0011111010;
    16'b0100010110000100: out_v[286] = 10'b0101011110;
    16'b0000100000010000: out_v[286] = 10'b1011101000;
    16'b1100110000000100: out_v[286] = 10'b1001000100;
    default: out_v[286] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000100000000001: out_v[287] = 10'b1001101110;
    16'b0010000000000001: out_v[287] = 10'b0011000001;
    16'b0000000000000001: out_v[287] = 10'b0011000001;
    16'b0100000000000001: out_v[287] = 10'b1100100111;
    16'b0010000000000000: out_v[287] = 10'b1110010011;
    16'b0100100000000001: out_v[287] = 10'b1000101001;
    16'b1010100000000001: out_v[287] = 10'b0010110011;
    16'b1100100100000001: out_v[287] = 10'b1101000010;
    16'b1000000000000001: out_v[287] = 10'b0100011011;
    16'b0000000000000000: out_v[287] = 10'b0010000101;
    16'b0000100000000000: out_v[287] = 10'b1001101100;
    16'b0110000000000001: out_v[287] = 10'b1100100110;
    16'b0010100000000001: out_v[287] = 10'b0000110110;
    16'b1010000000000001: out_v[287] = 10'b1000110111;
    16'b0100000000000000: out_v[287] = 10'b0010101010;
    16'b1000100000000001: out_v[287] = 10'b0111010111;
    16'b0100000100000001: out_v[287] = 10'b0111000011;
    16'b0100100100000001: out_v[287] = 10'b1000010011;
    16'b1100000100000001: out_v[287] = 10'b1001001000;
    16'b1100100100000000: out_v[287] = 10'b0010010110;
    16'b1000000100000001: out_v[287] = 10'b1000111111;
    16'b1000000000000000: out_v[287] = 10'b1010001111;
    16'b1000000100000000: out_v[287] = 10'b0100111010;
    16'b1100000100000000: out_v[287] = 10'b1011011010;
    16'b1000100100000001: out_v[287] = 10'b0111010000;
    16'b1000100000000000: out_v[287] = 10'b0011010110;
    16'b1110100100000000: out_v[287] = 10'b1000010111;
    16'b1000100100000000: out_v[287] = 10'b0111011000;
    16'b1100110100000001: out_v[287] = 10'b1110100100;
    16'b0100100100000000: out_v[287] = 10'b1000110010;
    16'b0010100000000000: out_v[287] = 10'b0000100111;
    16'b0100000100000000: out_v[287] = 10'b1011100110;
    16'b1100110100000000: out_v[287] = 10'b1001010100;
    16'b0100100000000000: out_v[287] = 10'b1000111011;
    16'b0000100100000001: out_v[287] = 10'b1100101100;
    16'b0100110100000000: out_v[287] = 10'b1110111011;
    16'b0100010100000000: out_v[287] = 10'b0011011101;
    16'b0000100100000000: out_v[287] = 10'b1000101110;
    16'b0110100100000001: out_v[287] = 10'b0110010001;
    16'b0010100100000001: out_v[287] = 10'b1100000110;
    16'b1110100100000001: out_v[287] = 10'b1110000100;
    16'b0100110100000001: out_v[287] = 10'b1001001110;
    16'b0010100100000000: out_v[287] = 10'b1110111011;
    16'b1110000100000000: out_v[287] = 10'b1101011000;
    16'b1100000000000001: out_v[287] = 10'b1001011101;
    16'b1110000100000001: out_v[287] = 10'b0011011100;
    16'b1100000000000000: out_v[287] = 10'b1111100100;
    16'b1100000100001000: out_v[287] = 10'b1001110011;
    16'b1100100000000001: out_v[287] = 10'b1111100100;
    16'b1100100000000000: out_v[287] = 10'b0111100011;
    16'b1010100100000000: out_v[287] = 10'b1100100100;
    16'b1010000100000001: out_v[287] = 10'b0011100100;
    16'b1010100100000001: out_v[287] = 10'b0011101000;
    16'b0110100100000000: out_v[287] = 10'b0100011111;
    16'b1010000100000000: out_v[287] = 10'b1100100010;
    16'b1010000000000000: out_v[287] = 10'b0101111101;
    16'b0000000100000001: out_v[287] = 10'b0111101000;
    16'b0000000100000000: out_v[287] = 10'b0101100000;
    16'b0110000100000001: out_v[287] = 10'b0010000011;
    16'b0010000100000001: out_v[287] = 10'b0011111110;
    default: out_v[287] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001100000001000: out_v[288] = 10'b0100100111;
    16'b0001001010001001: out_v[288] = 10'b0010001010;
    16'b0001001010101101: out_v[288] = 10'b1000101001;
    16'b0001101010101101: out_v[288] = 10'b0100100011;
    16'b0001001000001000: out_v[288] = 10'b1001011101;
    16'b0000100010001001: out_v[288] = 10'b0010100101;
    16'b0001001010001101: out_v[288] = 10'b1011000011;
    16'b0000001010101101: out_v[288] = 10'b0011001011;
    16'b0001100010001001: out_v[288] = 10'b0110001101;
    16'b0000001010001101: out_v[288] = 10'b0000011101;
    16'b0001101010001001: out_v[288] = 10'b1010111111;
    16'b0001001010000001: out_v[288] = 10'b0101010111;
    16'b0001101000001000: out_v[288] = 10'b0100110100;
    16'b0001101010001101: out_v[288] = 10'b0011000110;
    16'b0001000010001001: out_v[288] = 10'b1010100010;
    16'b0000000010001101: out_v[288] = 10'b1111100011;
    16'b0001000010001101: out_v[288] = 10'b1100101011;
    16'b0000000010001001: out_v[288] = 10'b1100111000;
    16'b0000001010001001: out_v[288] = 10'b1100100110;
    16'b0001101000001100: out_v[288] = 10'b0111011111;
    16'b0001000010101001: out_v[288] = 10'b0111000000;
    16'b0000000000001000: out_v[288] = 10'b0111011000;
    16'b0001001010101001: out_v[288] = 10'b1011100011;
    16'b0001100010001101: out_v[288] = 10'b1101000100;
    16'b0000101010001101: out_v[288] = 10'b0011100111;
    16'b0001000000001000: out_v[288] = 10'b0101010111;
    16'b0001001010000101: out_v[288] = 10'b0010110000;
    16'b0001000010101101: out_v[288] = 10'b0101100001;
    16'b0100000010001001: out_v[288] = 10'b1001100100;
    16'b0001001000001100: out_v[288] = 10'b1110111011;
    16'b0001000000000000: out_v[288] = 10'b0011000110;
    16'b0000000000000000: out_v[288] = 10'b0011010001;
    16'b0000000010001000: out_v[288] = 10'b0011111101;
    16'b0100100010001001: out_v[288] = 10'b1001011011;
    16'b0001100010000001: out_v[288] = 10'b0110100110;
    16'b0000101010001001: out_v[288] = 10'b1010000100;
    16'b0000100010000001: out_v[288] = 10'b1110001110;
    16'b0000001010000001: out_v[288] = 10'b1110100010;
    16'b0000000010000001: out_v[288] = 10'b1101001101;
    16'b0000001000001000: out_v[288] = 10'b1011000101;
    16'b0000001000000000: out_v[288] = 10'b0011001110;
    16'b0000000011001001: out_v[288] = 10'b0000111111;
    16'b0000101010000001: out_v[288] = 10'b0100010101;
    16'b0001000011001001: out_v[288] = 10'b1011010100;
    16'b0000101011001001: out_v[288] = 10'b1011100110;
    16'b0001100011001001: out_v[288] = 10'b1010111111;
    16'b0000100000001000: out_v[288] = 10'b1011001010;
    16'b0000101000001000: out_v[288] = 10'b0111000010;
    16'b0000100011001001: out_v[288] = 10'b1111100011;
    16'b0001001000000000: out_v[288] = 10'b0011001011;
    16'b0001100000000000: out_v[288] = 10'b0010101000;
    16'b0001000010001000: out_v[288] = 10'b0001000101;
    16'b0001101000000000: out_v[288] = 10'b0001011011;
    16'b0001000010000001: out_v[288] = 10'b0110010110;
    16'b0001001010001000: out_v[288] = 10'b1010110111;
    16'b0000100000000100: out_v[288] = 10'b1000111001;
    16'b0000001000000100: out_v[288] = 10'b0101011100;
    16'b0000100000000000: out_v[288] = 10'b1001101010;
    16'b0000000000000100: out_v[288] = 10'b1111100000;
    16'b0001100000000100: out_v[288] = 10'b0001110100;
    16'b0100100000001100: out_v[288] = 10'b0001111111;
    16'b0000101000100100: out_v[288] = 10'b1010100011;
    16'b0001000000000100: out_v[288] = 10'b1001101100;
    16'b0001100000100100: out_v[288] = 10'b1101110000;
    16'b0000000000100100: out_v[288] = 10'b1001011001;
    16'b0000100000001100: out_v[288] = 10'b0011111111;
    16'b0001000000100100: out_v[288] = 10'b1011001100;
    16'b0101100000000000: out_v[288] = 10'b0101000111;
    16'b0000101001100100: out_v[288] = 10'b1010001000;
    16'b0100100000001000: out_v[288] = 10'b0101010010;
    16'b0000100000100100: out_v[288] = 10'b0010001011;
    16'b0000101000000000: out_v[288] = 10'b0000010101;
    16'b0100100000000000: out_v[288] = 10'b1111010101;
    16'b0000101000000100: out_v[288] = 10'b1111000010;
    16'b0000101001100000: out_v[288] = 10'b1101100110;
    16'b0101100000000100: out_v[288] = 10'b1101101101;
    16'b0101100000100100: out_v[288] = 10'b0011001101;
    16'b1000000010001001: out_v[288] = 10'b1010111011;
    16'b0001001000000100: out_v[288] = 10'b0100110100;
    16'b0001000000001100: out_v[288] = 10'b1001101010;
    16'b0101001010001101: out_v[288] = 10'b1101100010;
    16'b0101000010001001: out_v[288] = 10'b1000110101;
    16'b0101000000001000: out_v[288] = 10'b1111100010;
    16'b0101000010001101: out_v[288] = 10'b1011111000;
    16'b1001000000000000: out_v[288] = 10'b1011010011;
    16'b1001000010001001: out_v[288] = 10'b1011111110;
    16'b1101000010001001: out_v[288] = 10'b1000101110;
    16'b0101000000000000: out_v[288] = 10'b0110110111;
    16'b1001000000000100: out_v[288] = 10'b0110011111;
    16'b0001001000100100: out_v[288] = 10'b0110100000;
    16'b0101001010101101: out_v[288] = 10'b1011001001;
    16'b0001001000101100: out_v[288] = 10'b1010001010;
    16'b0101001010001001: out_v[288] = 10'b0001101000;
    16'b1001000010001101: out_v[288] = 10'b1011111110;
    16'b0000001000001100: out_v[288] = 10'b1001111010;
    16'b0010001010001001: out_v[288] = 10'b1100110011;
    16'b0010000010001001: out_v[288] = 10'b0111011000;
    16'b0000001000100100: out_v[288] = 10'b1001010110;
    16'b0000101010101101: out_v[288] = 10'b0101011110;
    16'b0000001010001000: out_v[288] = 10'b0000110110;
    16'b0000101000001100: out_v[288] = 10'b0101010111;
    16'b0000100000101100: out_v[288] = 10'b1011111110;
    16'b0001101000100100: out_v[288] = 10'b1111010111;
    16'b0001100000101100: out_v[288] = 10'b1110001111;
    16'b0001000000100000: out_v[288] = 10'b1000110001;
    16'b0001100000100000: out_v[288] = 10'b0010110000;
    16'b0000000000001100: out_v[288] = 10'b1101111110;
    16'b0000100000100000: out_v[288] = 10'b1001000011;
    16'b0001100000001100: out_v[288] = 10'b0110100010;
    16'b0101100010001001: out_v[288] = 10'b0011001110;
    16'b0001100010101101: out_v[288] = 10'b0101010010;
    16'b0001101000101100: out_v[288] = 10'b1001010110;
    16'b0000001001100100: out_v[288] = 10'b1010110010;
    16'b0000000000100000: out_v[288] = 10'b1101010011;
    default: out_v[288] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1010000000110000: out_v[289] = 10'b1000110011;
    16'b0000000000110000: out_v[289] = 10'b1010100111;
    16'b1010001000010001: out_v[289] = 10'b0101100111;
    16'b0010000000000000: out_v[289] = 10'b1110001001;
    16'b0000100000110000: out_v[289] = 10'b0011110001;
    16'b1010000000010000: out_v[289] = 10'b1010011011;
    16'b0000000000010000: out_v[289] = 10'b1010001111;
    16'b1000001000011001: out_v[289] = 10'b0100011101;
    16'b0010000000100000: out_v[289] = 10'b1101001001;
    16'b0010000000110000: out_v[289] = 10'b0110011000;
    16'b0000000000100000: out_v[289] = 10'b0011110000;
    16'b1010001000111001: out_v[289] = 10'b1000001001;
    16'b1010001000101001: out_v[289] = 10'b1000101100;
    16'b1010001000110001: out_v[289] = 10'b1001010111;
    16'b1010000000100000: out_v[289] = 10'b0001110111;
    16'b1010001000011001: out_v[289] = 10'b0100000101;
    16'b1010000000110001: out_v[289] = 10'b0111010011;
    16'b0010000000010000: out_v[289] = 10'b1001001100;
    16'b0010001000010000: out_v[289] = 10'b0010110111;
    16'b1010001000010000: out_v[289] = 10'b0011001101;
    16'b0000100000100000: out_v[289] = 10'b0111000100;
    16'b0010100000110000: out_v[289] = 10'b0100011110;
    16'b1010001000100001: out_v[289] = 10'b1011010011;
    16'b0010001000110000: out_v[289] = 10'b0110111000;
    16'b1010000000100001: out_v[289] = 10'b0101110010;
    16'b1010001000000001: out_v[289] = 10'b0101100110;
    16'b1010001000110000: out_v[289] = 10'b0111001010;
    16'b0010001000011000: out_v[289] = 10'b1010100100;
    16'b1010001000001001: out_v[289] = 10'b1000001101;
    16'b0000000000000000: out_v[289] = 10'b0011110110;
    16'b1000000000000000: out_v[289] = 10'b0100010011;
    16'b1010000000000000: out_v[289] = 10'b1010000101;
    16'b1000000000000001: out_v[289] = 10'b0100011100;
    16'b1010000000000001: out_v[289] = 10'b0110111111;
    16'b0010001000000001: out_v[289] = 10'b0010001001;
    16'b0000100000010000: out_v[289] = 10'b1001111011;
    16'b1000000000010001: out_v[289] = 10'b0011011011;
    16'b1000001000001001: out_v[289] = 10'b1111100100;
    16'b0010001000000000: out_v[289] = 10'b1111000101;
    16'b1000000000010000: out_v[289] = 10'b0110110000;
    16'b1000001000000001: out_v[289] = 10'b1011001101;
    16'b1000000000001001: out_v[289] = 10'b1111110010;
    16'b1000001000010001: out_v[289] = 10'b0110011001;
    16'b0010001000001000: out_v[289] = 10'b0010100000;
    16'b1010000000010001: out_v[289] = 10'b0110100011;
    16'b1000001000101001: out_v[289] = 10'b1110001110;
    16'b0010001000001001: out_v[289] = 10'b0100111101;
    16'b1000001000100001: out_v[289] = 10'b0110001101;
    16'b0010001000101001: out_v[289] = 10'b0001011110;
    16'b0010001000101000: out_v[289] = 10'b1010101110;
    16'b1000001000111001: out_v[289] = 10'b1100001000;
    16'b0010001000111000: out_v[289] = 10'b0010110000;
    16'b1000000000100001: out_v[289] = 10'b1010001100;
    16'b0010001000100000: out_v[289] = 10'b1100111010;
    16'b1000000000101001: out_v[289] = 10'b1010101010;
    16'b1000000000110001: out_v[289] = 10'b0001101010;
    16'b0000000000101000: out_v[289] = 10'b0001010010;
    16'b0000000000001000: out_v[289] = 10'b0011010011;
    16'b0000000000011000: out_v[289] = 10'b0101010010;
    16'b0000001000101000: out_v[289] = 10'b0101010000;
    16'b0000000000111000: out_v[289] = 10'b1001010000;
    16'b0000001000011000: out_v[289] = 10'b0011111100;
    16'b0000001000001000: out_v[289] = 10'b0000011011;
    16'b0000001000111000: out_v[289] = 10'b1001110011;
    16'b0010001000100001: out_v[289] = 10'b0001011000;
    16'b0000001000100000: out_v[289] = 10'b0111011011;
    16'b0010001000110001: out_v[289] = 10'b0001110110;
    16'b0010100000010000: out_v[289] = 10'b0111011100;
    16'b1010101000100001: out_v[289] = 10'b0000001010;
    16'b0010100000100000: out_v[289] = 10'b0111001011;
    16'b1010101000110001: out_v[289] = 10'b1111001101;
    16'b0010101000100000: out_v[289] = 10'b0111111111;
    16'b0010101000110000: out_v[289] = 10'b1101001011;
    16'b1010101000101001: out_v[289] = 10'b1011111111;
    16'b0000100000000000: out_v[289] = 10'b1000110101;
    16'b1010100000100000: out_v[289] = 10'b1010100100;
    16'b1010001000100000: out_v[289] = 10'b1000101101;
    16'b0011000000100000: out_v[289] = 10'b1111001010;
    16'b1011000000100000: out_v[289] = 10'b1011101010;
    16'b1011001000000001: out_v[289] = 10'b1110111011;
    16'b1011001000100001: out_v[289] = 10'b0111001111;
    16'b1011000000100001: out_v[289] = 10'b1111001101;
    16'b0001000000100000: out_v[289] = 10'b1101110100;
    16'b0000001000101001: out_v[289] = 10'b0011001011;
    16'b0001000000000000: out_v[289] = 10'b0011000111;
    16'b0000001000001001: out_v[289] = 10'b1011110010;
    16'b0010000010010000: out_v[289] = 10'b1111011011;
    16'b0010000000001000: out_v[289] = 10'b1111100001;
    16'b0010000010010010: out_v[289] = 10'b0000011111;
    16'b0000000010010000: out_v[289] = 10'b1111111011;
    16'b1010001000000000: out_v[289] = 10'b0010001100;
    default: out_v[289] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000010000010: out_v[290] = 10'b0101000111;
    16'b0000100000001011: out_v[290] = 10'b0001011011;
    16'b0000100010001011: out_v[290] = 10'b0111010011;
    16'b0000100000011011: out_v[290] = 10'b1111011001;
    16'b0000000010011010: out_v[290] = 10'b1011001101;
    16'b0000000010001010: out_v[290] = 10'b1010110101;
    16'b0000100010000011: out_v[290] = 10'b0110010101;
    16'b0000100010001111: out_v[290] = 10'b1011011100;
    16'b0000100000011001: out_v[290] = 10'b0100100011;
    16'b0000100000000010: out_v[290] = 10'b1101100101;
    16'b0000000010010110: out_v[290] = 10'b0100110101;
    16'b0000100010001001: out_v[290] = 10'b1110001111;
    16'b0000100010011111: out_v[290] = 10'b1101100111;
    16'b0000100000001010: out_v[290] = 10'b1001010101;
    16'b0000100000001000: out_v[290] = 10'b0110100111;
    16'b0000000000000010: out_v[290] = 10'b1001011001;
    16'b0000100000000011: out_v[290] = 10'b0101010011;
    16'b0000000000000011: out_v[290] = 10'b1100000111;
    16'b0000000010000011: out_v[290] = 10'b0000110001;
    16'b0000100010011011: out_v[290] = 10'b0110001001;
    16'b0000000000001000: out_v[290] = 10'b0010111100;
    16'b0000100010000010: out_v[290] = 10'b1100011001;
    16'b0000000010010010: out_v[290] = 10'b1100000101;
    16'b0000100010010011: out_v[290] = 10'b1110011111;
    16'b0000100000010011: out_v[290] = 10'b1111110111;
    16'b0000100010001110: out_v[290] = 10'b0011110110;
    16'b0000000000010010: out_v[290] = 10'b0110001011;
    16'b0000000010001110: out_v[290] = 10'b1111010010;
    16'b0000000000010011: out_v[290] = 10'b0010011011;
    16'b0000000000011000: out_v[290] = 10'b1001110111;
    16'b0000100000001001: out_v[290] = 10'b1001000001;
    16'b0000000010010011: out_v[290] = 10'b0110110010;
    16'b0000000000001010: out_v[290] = 10'b0001111000;
    16'b0000100000011010: out_v[290] = 10'b1111011101;
    16'b0000100000001111: out_v[290] = 10'b0000110110;
    16'b0000100010001010: out_v[290] = 10'b0011110000;
    16'b0000100000001110: out_v[290] = 10'b0110010100;
    16'b0000000000011010: out_v[290] = 10'b0011100101;
    16'b0000100010000111: out_v[290] = 10'b1100100111;
    16'b0000000010011110: out_v[290] = 10'b1111000001;
    16'b0000100010011001: out_v[290] = 10'b1110001011;
    16'b0000000000001110: out_v[290] = 10'b0000111110;
    16'b0000000010000110: out_v[290] = 10'b1110010010;
    16'b0000000000000000: out_v[290] = 10'b0111011100;
    16'b0000000000010000: out_v[290] = 10'b0110110010;
    16'b0000000010000000: out_v[290] = 10'b0101010100;
    16'b0000000000010100: out_v[290] = 10'b0010110000;
    16'b0000000000000100: out_v[290] = 10'b1010010010;
    16'b0000000010000100: out_v[290] = 10'b0101010100;
    16'b0000000010010000: out_v[290] = 10'b1000110010;
    16'b0000000010010100: out_v[290] = 10'b1001101001;
    16'b0010100010010110: out_v[290] = 10'b0011011110;
    16'b0010000010010010: out_v[290] = 10'b1100010100;
    16'b0010000010000000: out_v[290] = 10'b1010100101;
    16'b0000100010010110: out_v[290] = 10'b1001111001;
    16'b0000000000010110: out_v[290] = 10'b0011001111;
    16'b0000100010011100: out_v[290] = 10'b1010101010;
    16'b0000100010011110: out_v[290] = 10'b1011011010;
    16'b0010000010010110: out_v[290] = 10'b1110011101;
    16'b0000000010011100: out_v[290] = 10'b1111000111;
    16'b0000100010011010: out_v[290] = 10'b0010001110;
    16'b0000100010000110: out_v[290] = 10'b1001101100;
    16'b0000100010000100: out_v[290] = 10'b0101111000;
    16'b0000000000000110: out_v[290] = 10'b1011101011;
    16'b0000100000010110: out_v[290] = 10'b0010001100;
    16'b0000100000011100: out_v[290] = 10'b0110100110;
    16'b0000100010011101: out_v[290] = 10'b1010110101;
    16'b0010000010010000: out_v[290] = 10'b1011100010;
    16'b0010000010000100: out_v[290] = 10'b0010100111;
    16'b0000100010001100: out_v[290] = 10'b0010111111;
    16'b0010000010000010: out_v[290] = 10'b1111010110;
    16'b0000100010010111: out_v[290] = 10'b0110000101;
    16'b0000100010010010: out_v[290] = 10'b1010011100;
    16'b0000000000100000: out_v[290] = 10'b1111001101;
    16'b0000001000000110: out_v[290] = 10'b1011110010;
    16'b0000001000000010: out_v[290] = 10'b0000110010;
    16'b0000000010100000: out_v[290] = 10'b1100001000;
    16'b0000000000011110: out_v[290] = 10'b1111011011;
    16'b0000100000010010: out_v[290] = 10'b0001001110;
    16'b0000001000001110: out_v[290] = 10'b1011011011;
    16'b0000000000100010: out_v[290] = 10'b0011001110;
    16'b0000000000100110: out_v[290] = 10'b1111100101;
    16'b0000001000000100: out_v[290] = 10'b1011001000;
    16'b0000100000011110: out_v[290] = 10'b1100111000;
    16'b0000000000001100: out_v[290] = 10'b1001101001;
    16'b0000000000100100: out_v[290] = 10'b0001010101;
    16'b0000000000000101: out_v[290] = 10'b0100011111;
    16'b0000000000001111: out_v[290] = 10'b0000100010;
    16'b0000001000000101: out_v[290] = 10'b0001111111;
    16'b0000000010000101: out_v[290] = 10'b0101000111;
    16'b0000000000000111: out_v[290] = 10'b0001111100;
    16'b0000000010001111: out_v[290] = 10'b0110010110;
    16'b0000000000001101: out_v[290] = 10'b0101100000;
    16'b0000100000001101: out_v[290] = 10'b1001011011;
    16'b0000100000000111: out_v[290] = 10'b0111110110;
    16'b0000100000000101: out_v[290] = 10'b1001101011;
    16'b0000000010001101: out_v[290] = 10'b0110110011;
    16'b0000000010001100: out_v[290] = 10'b1100001100;
    16'b0000001000001111: out_v[290] = 10'b1011100111;
    16'b0000100010000101: out_v[290] = 10'b0101110010;
    16'b0000100000000110: out_v[290] = 10'b1111001010;
    16'b0000001000001010: out_v[290] = 10'b0011110000;
    16'b0000100010000000: out_v[290] = 10'b1101111011;
    16'b0000000000011100: out_v[290] = 10'b1111010010;
    16'b0000000000001011: out_v[290] = 10'b0000101000;
    16'b0000100000011000: out_v[290] = 10'b0110110001;
    16'b0000100010010101: out_v[290] = 10'b0001011000;
    16'b0000000010010001: out_v[290] = 10'b0011000000;
    16'b0000000010000001: out_v[290] = 10'b1101000101;
    16'b0000100010010001: out_v[290] = 10'b0011110010;
    16'b0000000010010101: out_v[290] = 10'b1110111111;
    16'b0000100010010100: out_v[290] = 10'b0011011010;
    16'b0000100010000001: out_v[290] = 10'b1011011011;
    16'b0000000011000110: out_v[290] = 10'b0011000001;
    16'b0000001000100110: out_v[290] = 10'b0000011110;
    16'b0000000001000110: out_v[290] = 10'b1100000101;
    16'b0000001010000110: out_v[290] = 10'b1010100010;
    16'b0000001000000111: out_v[290] = 10'b1001001000;
    16'b0000001000000000: out_v[290] = 10'b0001001111;
    16'b0000001010001110: out_v[290] = 10'b0111010001;
    16'b0000000010001000: out_v[290] = 10'b1010100011;
    16'b0000100000001100: out_v[290] = 10'b0101010101;
    16'b0000000000000001: out_v[290] = 10'b1010101110;
    16'b0000000010000111: out_v[290] = 10'b1001111011;
    default: out_v[290] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100000010010001: out_v[291] = 10'b1101000101;
    16'b1100000010010000: out_v[291] = 10'b1110000110;
    16'b1100000110010010: out_v[291] = 10'b0010011010;
    16'b0000000010010000: out_v[291] = 10'b0000011001;
    16'b1100100010010010: out_v[291] = 10'b1100010110;
    16'b1100000010010010: out_v[291] = 10'b1100010001;
    16'b0100000010000000: out_v[291] = 10'b0000100101;
    16'b1000000010000000: out_v[291] = 10'b1101101001;
    16'b0100100010000000: out_v[291] = 10'b1011100011;
    16'b1100000000000010: out_v[291] = 10'b0000001011;
    16'b1100000010000000: out_v[291] = 10'b1011110010;
    16'b1100000010010011: out_v[291] = 10'b1001001111;
    16'b0100000000000000: out_v[291] = 10'b1110100000;
    16'b0100000010010000: out_v[291] = 10'b1110001001;
    16'b0100100010010000: out_v[291] = 10'b0110000111;
    16'b0100000010010010: out_v[291] = 10'b1000111011;
    16'b1000000010010000: out_v[291] = 10'b0001011100;
    16'b1100100110010010: out_v[291] = 10'b1100011111;
    16'b1100000000000000: out_v[291] = 10'b0010100111;
    16'b1100100010010000: out_v[291] = 10'b1100000111;
    16'b1100000000010010: out_v[291] = 10'b1000011000;
    16'b0100100100010000: out_v[291] = 10'b1000001001;
    16'b0100100010010010: out_v[291] = 10'b1010001111;
    16'b0100000000010000: out_v[291] = 10'b1111011101;
    16'b1100000000010001: out_v[291] = 10'b0001011101;
    16'b1100100110010000: out_v[291] = 10'b0010011111;
    16'b0100100100000000: out_v[291] = 10'b0011100001;
    16'b0000000010000000: out_v[291] = 10'b1000010110;
    16'b0100000010000010: out_v[291] = 10'b0010011000;
    16'b1100000010000010: out_v[291] = 10'b0011011100;
    16'b1100000000010000: out_v[291] = 10'b1110001001;
    16'b1100000000010011: out_v[291] = 10'b0100010111;
    16'b1100000110010000: out_v[291] = 10'b0001101110;
    16'b1100000010010001: out_v[291] = 10'b1101100011;
    16'b1100000000000011: out_v[291] = 10'b0001110111;
    16'b0100000000010011: out_v[291] = 10'b0011010010;
    16'b0100000000010010: out_v[291] = 10'b1000011111;
    16'b1000000000000000: out_v[291] = 10'b0110100110;
    16'b0100000000000010: out_v[291] = 10'b0110001001;
    16'b0000000000000011: out_v[291] = 10'b0100100100;
    16'b0000000000010010: out_v[291] = 10'b0011101010;
    16'b1000000000000010: out_v[291] = 10'b1100110010;
    16'b0000000000000000: out_v[291] = 10'b0000101110;
    16'b0100000000000011: out_v[291] = 10'b1110011000;
    16'b0000000000010011: out_v[291] = 10'b0000110010;
    16'b0000000000000010: out_v[291] = 10'b0001111101;
    16'b1100100000010000: out_v[291] = 10'b0011010100;
    16'b1100100000000010: out_v[291] = 10'b0111110010;
    16'b1000000000010000: out_v[291] = 10'b0001011111;
    16'b1100100000000011: out_v[291] = 10'b1001111100;
    16'b1100100000010001: out_v[291] = 10'b1111011001;
    16'b1000000000010001: out_v[291] = 10'b0110111100;
    16'b1100100000010011: out_v[291] = 10'b1000000111;
    16'b1000100000010000: out_v[291] = 10'b0101010101;
    16'b0100100000010011: out_v[291] = 10'b1011111111;
    16'b0100000000010001: out_v[291] = 10'b1110001101;
    16'b1000100000010001: out_v[291] = 10'b0111011111;
    16'b0100100000000010: out_v[291] = 10'b1010001100;
    16'b0100100000010001: out_v[291] = 10'b0111011011;
    16'b0000100000010000: out_v[291] = 10'b1101011110;
    16'b1100100000010010: out_v[291] = 10'b1011001010;
    16'b1000000000000001: out_v[291] = 10'b0001001110;
    16'b0000000000010000: out_v[291] = 10'b0001011110;
    16'b1100000000000001: out_v[291] = 10'b1111101000;
    16'b0000000000010001: out_v[291] = 10'b0100111011;
    16'b0000100000010001: out_v[291] = 10'b1100111000;
    16'b0100000000000001: out_v[291] = 10'b1101100110;
    16'b0100100000010000: out_v[291] = 10'b1100000110;
    16'b0100100000000011: out_v[291] = 10'b0111001011;
    16'b0000000000000001: out_v[291] = 10'b0011011111;
    16'b1000100000000011: out_v[291] = 10'b1100110110;
    16'b0100000000001010: out_v[291] = 10'b0000000011;
    16'b0100100010000010: out_v[291] = 10'b1111011011;
    16'b1000000000010010: out_v[291] = 10'b1011001011;
    16'b0100100000010010: out_v[291] = 10'b1011011010;
    16'b0100000010010011: out_v[291] = 10'b1101000000;
    16'b0100000010000011: out_v[291] = 10'b0001011111;
    16'b1100000010000011: out_v[291] = 10'b0100111101;
    16'b1000000010011000: out_v[291] = 10'b0001111011;
    16'b1000000010000010: out_v[291] = 10'b1101110010;
    16'b0000000010010011: out_v[291] = 10'b1100100111;
    16'b1000000010010001: out_v[291] = 10'b0110001101;
    16'b0000000010010001: out_v[291] = 10'b0100111111;
    16'b0000000010010010: out_v[291] = 10'b0110100111;
    16'b1000000000000011: out_v[291] = 10'b0101010000;
    16'b0000000010000001: out_v[291] = 10'b1111010110;
    16'b0000100100010001: out_v[291] = 10'b0110110011;
    16'b1000000010010010: out_v[291] = 10'b1011101000;
    16'b0000000010000010: out_v[291] = 10'b1100100101;
    16'b0000000010000011: out_v[291] = 10'b1000101011;
    16'b0000000100010000: out_v[291] = 10'b1011001011;
    16'b0000000100010001: out_v[291] = 10'b0100111101;
    16'b1000000010010011: out_v[291] = 10'b1001100010;
    16'b1000000010011001: out_v[291] = 10'b0101111110;
    16'b1000000010000011: out_v[291] = 10'b1001010110;
    16'b1000000010000001: out_v[291] = 10'b0011001011;
    16'b1100000010000001: out_v[291] = 10'b0000101100;
    16'b0100000010001001: out_v[291] = 10'b0000100110;
    16'b0100000010000001: out_v[291] = 10'b1010101010;
    16'b0000100010000000: out_v[291] = 10'b0111111010;
    16'b1000000000010011: out_v[291] = 10'b1111100001;
    16'b0100000010001000: out_v[291] = 10'b0000100110;
    16'b1000100010000001: out_v[291] = 10'b0011001011;
    16'b1000100010000000: out_v[291] = 10'b0110001001;
    16'b1100100010000001: out_v[291] = 10'b1011000000;
    16'b1100000010011010: out_v[291] = 10'b0011100010;
    16'b1000000010011010: out_v[291] = 10'b0011001110;
    16'b1100000000011010: out_v[291] = 10'b1110100000;
    16'b1000000000011010: out_v[291] = 10'b0011110011;
    16'b0000000110010010: out_v[291] = 10'b0011100100;
    16'b1100000100010000: out_v[291] = 10'b0000110101;
    16'b1000000110011010: out_v[291] = 10'b0111010101;
    16'b1100000000001010: out_v[291] = 10'b0011100000;
    16'b1100000000011000: out_v[291] = 10'b0010101010;
    16'b1100000110011010: out_v[291] = 10'b0010110000;
    16'b1000000000001010: out_v[291] = 10'b0011101001;
    16'b1100000100011000: out_v[291] = 10'b1010100011;
    16'b1100000000001011: out_v[291] = 10'b0011110100;
    16'b1100000100011010: out_v[291] = 10'b1101010010;
    16'b1000000100011010: out_v[291] = 10'b1111101011;
    16'b0000000110011010: out_v[291] = 10'b0001011011;
    16'b1100000010001010: out_v[291] = 10'b0111111111;
    16'b1100000010011000: out_v[291] = 10'b1011001010;
    16'b0100000110010010: out_v[291] = 10'b1111001011;
    16'b1000000110010010: out_v[291] = 10'b0100101110;
    16'b0000000010011010: out_v[291] = 10'b1110001100;
    16'b0000000100010010: out_v[291] = 10'b0111111101;
    16'b0100000010011000: out_v[291] = 10'b1101001110;
    16'b1100000010011001: out_v[291] = 10'b1101000111;
    16'b1100000010011011: out_v[291] = 10'b1101001010;
    16'b1100000010001001: out_v[291] = 10'b1101001101;
    16'b0100000100010011: out_v[291] = 10'b1100010111;
    16'b1100000000011001: out_v[291] = 10'b1101000101;
    16'b1100000010001011: out_v[291] = 10'b1101000011;
    16'b0100000100010001: out_v[291] = 10'b1101000101;
    16'b0100000010011001: out_v[291] = 10'b0001111000;
    16'b1100000010001000: out_v[291] = 10'b1100000010;
    default: out_v[291] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001000000010100: out_v[292] = 10'b0010100101;
    16'b0001000000011100: out_v[292] = 10'b1000110001;
    16'b0001000000011000: out_v[292] = 10'b0010000111;
    16'b0000000000001100: out_v[292] = 10'b0000110101;
    16'b0000000000000100: out_v[292] = 10'b0001001101;
    16'b0001001000011100: out_v[292] = 10'b1011100011;
    16'b0001101000011100: out_v[292] = 10'b0101010110;
    16'b0001000000001000: out_v[292] = 10'b1010110101;
    16'b0001000000001100: out_v[292] = 10'b1001111111;
    16'b0001100000010100: out_v[292] = 10'b1001000101;
    16'b0001000000000100: out_v[292] = 10'b0010111100;
    16'b0001000000010000: out_v[292] = 10'b0010110111;
    16'b0000000000011100: out_v[292] = 10'b1000110111;
    16'b0000100000010100: out_v[292] = 10'b1100101001;
    16'b0000000000010100: out_v[292] = 10'b0001001101;
    16'b0001000000000000: out_v[292] = 10'b1011001001;
    16'b0000000000000000: out_v[292] = 10'b1010101011;
    16'b0000000000001000: out_v[292] = 10'b1010110000;
    16'b0001100000011100: out_v[292] = 10'b0001001101;
    16'b0000101000000100: out_v[292] = 10'b0011111110;
    16'b0000001000000000: out_v[292] = 10'b1001000010;
    16'b0000001000000100: out_v[292] = 10'b1110100010;
    16'b0001001000010000: out_v[292] = 10'b1101111100;
    16'b0001101000010000: out_v[292] = 10'b0000110010;
    16'b0001001000010100: out_v[292] = 10'b0110010001;
    16'b0000101000000000: out_v[292] = 10'b0010011100;
    16'b0001001000000000: out_v[292] = 10'b1101001100;
    16'b0001101000010100: out_v[292] = 10'b1100000110;
    16'b0000101000010100: out_v[292] = 10'b1100001011;
    16'b0000001000010100: out_v[292] = 10'b1111000100;
    16'b0000101000001100: out_v[292] = 10'b1011000100;
    16'b0000100000000000: out_v[292] = 10'b1100011001;
    16'b0000101000001000: out_v[292] = 10'b1101010100;
    16'b0001101000000100: out_v[292] = 10'b0010100010;
    16'b0000100000000100: out_v[292] = 10'b1000001000;
    16'b0001100000011000: out_v[292] = 10'b0110111010;
    16'b0000100000001100: out_v[292] = 10'b1101100000;
    16'b0001101000001000: out_v[292] = 10'b0111101101;
    16'b0001101000000000: out_v[292] = 10'b1000101000;
    16'b0001001000000100: out_v[292] = 10'b0110110011;
    16'b0001101000001100: out_v[292] = 10'b0010101110;
    16'b0000001000001100: out_v[292] = 10'b0001001000;
    16'b0001001000011000: out_v[292] = 10'b0101110010;
    16'b0000001000001000: out_v[292] = 10'b0011111000;
    16'b0001100000000100: out_v[292] = 10'b0111011110;
    16'b0001101000011000: out_v[292] = 10'b1101000000;
    16'b0001100000010000: out_v[292] = 10'b0100010001;
    16'b0001001000001100: out_v[292] = 10'b0111110010;
    16'b0001100000001100: out_v[292] = 10'b0101101010;
    16'b0001001000001000: out_v[292] = 10'b1100011100;
    16'b0000101000011100: out_v[292] = 10'b1010011010;
    16'b0001111000011100: out_v[292] = 10'b0010111011;
    16'b0000100000001000: out_v[292] = 10'b0111001000;
    16'b0000101001000000: out_v[292] = 10'b0001011000;
    16'b0000101000010000: out_v[292] = 10'b0100111110;
    16'b0000000000010000: out_v[292] = 10'b0001101011;
    16'b0000100000011100: out_v[292] = 10'b0001010010;
    16'b0000001000011100: out_v[292] = 10'b1101011110;
    16'b0001000001011000: out_v[292] = 10'b0111100110;
    16'b0001111000010000: out_v[292] = 10'b0011001011;
    16'b0001101010010100: out_v[292] = 10'b0100110111;
    16'b0001110000010000: out_v[292] = 10'b1111101010;
    16'b0001111001010000: out_v[292] = 10'b1111111100;
    16'b0001010000010000: out_v[292] = 10'b1011111011;
    16'b0001110000010100: out_v[292] = 10'b1101011011;
    16'b0001111000010100: out_v[292] = 10'b1100101100;
    16'b0001101001010000: out_v[292] = 10'b1010001011;
    16'b0001110001010000: out_v[292] = 10'b0101001011;
    16'b0001100010010100: out_v[292] = 10'b0111101010;
    16'b0001010000011000: out_v[292] = 10'b0111000011;
    16'b0001000001010000: out_v[292] = 10'b0000111010;
    16'b0000100000010000: out_v[292] = 10'b0001001111;
    16'b0001010001011000: out_v[292] = 10'b0011111010;
    16'b0001101001000000: out_v[292] = 10'b1100000101;
    16'b0001100000000000: out_v[292] = 10'b1100011100;
    16'b0001101001011000: out_v[292] = 10'b1001100111;
    16'b0001100001010000: out_v[292] = 10'b0011111011;
    16'b0001100001000000: out_v[292] = 10'b1101111101;
    16'b0001001001010000: out_v[292] = 10'b1101100101;
    default: out_v[292] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1101001110100000: out_v[293] = 10'b1101110110;
    16'b1000000110100000: out_v[293] = 10'b1000010001;
    16'b1100001110101001: out_v[293] = 10'b0100101100;
    16'b0000001100100000: out_v[293] = 10'b0001000101;
    16'b1000000110000000: out_v[293] = 10'b1011111100;
    16'b1100001110001001: out_v[293] = 10'b1010101100;
    16'b1000000110001001: out_v[293] = 10'b0011010011;
    16'b1000000110001000: out_v[293] = 10'b1100011100;
    16'b1000001110101000: out_v[293] = 10'b0100110100;
    16'b1001001110100000: out_v[293] = 10'b0011110111;
    16'b1101001110101000: out_v[293] = 10'b0010110111;
    16'b1000001110100000: out_v[293] = 10'b1110011010;
    16'b1101001010101000: out_v[293] = 10'b1000010101;
    16'b0000001100101000: out_v[293] = 10'b0101011001;
    16'b1101001110101001: out_v[293] = 10'b0000000011;
    16'b1100001110001000: out_v[293] = 10'b1010011011;
    16'b1000001110001001: out_v[293] = 10'b1110110011;
    16'b1101001010101001: out_v[293] = 10'b1111010101;
    16'b1000000110101000: out_v[293] = 10'b1110010101;
    16'b1000100110000000: out_v[293] = 10'b1100110010;
    16'b1100001110101000: out_v[293] = 10'b1001111110;
    16'b1100000110101000: out_v[293] = 10'b0010010101;
    16'b1000100110100000: out_v[293] = 10'b0010011001;
    16'b1101001000101000: out_v[293] = 10'b1010101110;
    16'b1000100110001000: out_v[293] = 10'b0111010111;
    16'b1100000110001001: out_v[293] = 10'b0010101111;
    16'b1101001100101000: out_v[293] = 10'b1011111111;
    16'b0100001100101000: out_v[293] = 10'b1101111110;
    16'b1101001010100000: out_v[293] = 10'b0011010011;
    16'b1000001110001000: out_v[293] = 10'b1100011010;
    16'b1101000010101000: out_v[293] = 10'b1011011011;
    16'b1100001010101001: out_v[293] = 10'b1011110100;
    16'b1100001110100000: out_v[293] = 10'b1111011100;
    16'b0000000000010000: out_v[293] = 10'b0010000111;
    16'b1000000010110000: out_v[293] = 10'b0101010100;
    16'b1001000010110000: out_v[293] = 10'b0011001110;
    16'b1001000010010000: out_v[293] = 10'b1000110111;
    16'b1001101110010000: out_v[293] = 10'b1011000010;
    16'b0001001010010000: out_v[293] = 10'b1111110011;
    16'b1001001010110000: out_v[293] = 10'b1001111110;
    16'b1000000000010000: out_v[293] = 10'b0100001010;
    16'b1000100010110000: out_v[293] = 10'b1010000010;
    16'b1000000010010000: out_v[293] = 10'b1100110001;
    16'b0000000010010000: out_v[293] = 10'b0010110101;
    16'b1001100110110000: out_v[293] = 10'b0101010001;
    16'b0000000010110000: out_v[293] = 10'b0111010000;
    16'b0001000010010000: out_v[293] = 10'b0011001101;
    16'b1000000000110000: out_v[293] = 10'b0001011011;
    16'b0000000000110000: out_v[293] = 10'b0000010111;
    16'b0001101110010000: out_v[293] = 10'b0011010011;
    16'b1001101110110000: out_v[293] = 10'b0011111111;
    16'b0001001010110000: out_v[293] = 10'b1001000111;
    16'b1000001010110000: out_v[293] = 10'b0111100000;
    16'b1001100010110000: out_v[293] = 10'b0011100110;
    16'b1100000110010000: out_v[293] = 10'b0000101101;
    16'b0000000100010000: out_v[293] = 10'b1001000011;
    16'b1100001100010000: out_v[293] = 10'b1011101011;
    16'b0000100000010000: out_v[293] = 10'b1001100101;
    16'b1100100110010000: out_v[293] = 10'b0010010111;
    16'b0100000100010000: out_v[293] = 10'b0100001011;
    16'b1000100100010000: out_v[293] = 10'b0010110001;
    16'b1100001110010000: out_v[293] = 10'b1000101110;
    16'b0100100100010000: out_v[293] = 10'b1110000111;
    16'b0001000000110000: out_v[293] = 10'b1111100100;
    16'b0000100000000000: out_v[293] = 10'b0110001101;
    16'b0100101100010000: out_v[293] = 10'b0011100101;
    16'b1100101110000000: out_v[293] = 10'b0011110100;
    16'b1100101110010000: out_v[293] = 10'b0101001101;
    16'b0000100100000000: out_v[293] = 10'b1101001110;
    16'b0100100100000000: out_v[293] = 10'b1100111011;
    16'b1000100010000000: out_v[293] = 10'b0111011101;
    16'b1000100010010000: out_v[293] = 10'b1001101101;
    16'b1100101100000000: out_v[293] = 10'b1111010001;
    16'b1100001110110000: out_v[293] = 10'b0010111000;
    16'b1000100100000000: out_v[293] = 10'b1110110011;
    16'b0100000100000000: out_v[293] = 10'b1101100110;
    16'b1000100000010000: out_v[293] = 10'b0111000100;
    16'b1100000100010000: out_v[293] = 10'b1011100001;
    16'b1000101010010000: out_v[293] = 10'b1010001001;
    16'b1000101110010000: out_v[293] = 10'b1110001010;
    16'b1000100110010000: out_v[293] = 10'b0110110101;
    16'b1100101100010000: out_v[293] = 10'b1010110111;
    16'b0000101100000000: out_v[293] = 10'b0011110010;
    16'b0100001100010000: out_v[293] = 10'b1111010110;
    16'b1100100100000000: out_v[293] = 10'b1111100111;
    16'b1100101110110000: out_v[293] = 10'b1110110101;
    16'b1000101010000000: out_v[293] = 10'b0100101110;
    16'b0000100100010000: out_v[293] = 10'b1001010101;
    16'b1000101110000000: out_v[293] = 10'b1101000111;
    16'b1100100100010000: out_v[293] = 10'b1010111011;
    16'b1000001110010000: out_v[293] = 10'b1100011011;
    16'b1100100110000000: out_v[293] = 10'b0111011001;
    16'b0100101100000000: out_v[293] = 10'b1001000001;
    16'b0000000100000000: out_v[293] = 10'b1110001110;
    16'b0000101000010000: out_v[293] = 10'b0001101111;
    16'b0100000000010000: out_v[293] = 10'b1001111100;
    16'b1101001100110000: out_v[293] = 10'b1001011000;
    16'b1000100100110000: out_v[293] = 10'b0111010010;
    16'b1001001110110000: out_v[293] = 10'b0100111110;
    16'b1101001110110000: out_v[293] = 10'b0010111110;
    16'b0100000100110000: out_v[293] = 10'b1111010101;
    16'b1101101110110000: out_v[293] = 10'b0101011001;
    16'b1101001010110000: out_v[293] = 10'b0010100111;
    16'b0101000000110000: out_v[293] = 10'b1001101011;
    16'b0000000100100000: out_v[293] = 10'b1011000111;
    16'b1000101110110000: out_v[293] = 10'b0100001000;
    16'b1101000110110000: out_v[293] = 10'b1111010011;
    16'b1101000110100000: out_v[293] = 10'b1001011110;
    16'b0000001100110000: out_v[293] = 10'b1100100011;
    16'b0000100100110000: out_v[293] = 10'b1011000101;
    16'b1000100110110000: out_v[293] = 10'b0110011000;
    16'b1001001100110000: out_v[293] = 10'b0010111101;
    16'b1101000000110000: out_v[293] = 10'b0111100011;
    16'b1000101100110000: out_v[293] = 10'b1100100111;
    16'b1101001000110000: out_v[293] = 10'b0000110010;
    16'b1000000110110000: out_v[293] = 10'b0010001110;
    16'b1000000100110000: out_v[293] = 10'b1110110101;
    16'b1101000100110000: out_v[293] = 10'b0111110000;
    16'b1101000010110000: out_v[293] = 10'b1110011001;
    16'b0101000100110000: out_v[293] = 10'b0011111111;
    16'b1100001100110000: out_v[293] = 10'b0000101110;
    16'b1000001110110000: out_v[293] = 10'b0001011101;
    16'b1000001100110000: out_v[293] = 10'b1111010010;
    16'b1101101010110000: out_v[293] = 10'b0010111011;
    16'b0000101100110000: out_v[293] = 10'b0101011010;
    16'b1101000010100000: out_v[293] = 10'b0111011110;
    16'b1001100100110000: out_v[293] = 10'b0001111110;
    16'b0000000100110000: out_v[293] = 10'b0010101111;
    16'b1001101100110000: out_v[293] = 10'b0111010010;
    16'b1100000110110000: out_v[293] = 10'b1111010111;
    16'b1101001110111000: out_v[293] = 10'b1010011110;
    16'b1101100100110000: out_v[293] = 10'b1011011011;
    16'b1000000110010000: out_v[293] = 10'b0001001010;
    16'b1101101100110000: out_v[293] = 10'b0111011011;
    16'b0100000100100000: out_v[293] = 10'b0011100100;
    16'b0000100100011000: out_v[293] = 10'b1110101111;
    16'b0000100000111001: out_v[293] = 10'b0101011111;
    16'b0000101000111000: out_v[293] = 10'b0001111101;
    16'b0000000100011000: out_v[293] = 10'b0111110111;
    16'b0100100100001000: out_v[293] = 10'b1011011001;
    16'b0000101000110000: out_v[293] = 10'b0100010101;
    16'b0000100000011000: out_v[293] = 10'b1000110100;
    16'b0001100100111000: out_v[293] = 10'b0101110011;
    16'b0001100100011001: out_v[293] = 10'b1111001101;
    16'b0000100000110000: out_v[293] = 10'b0010110001;
    16'b0000100010110000: out_v[293] = 10'b0010111101;
    16'b0000100000111000: out_v[293] = 10'b0111110000;
    16'b0000100010011000: out_v[293] = 10'b0111101101;
    16'b0001100100011000: out_v[293] = 10'b0010101001;
    16'b0100100100011000: out_v[293] = 10'b0100010111;
    16'b0001100000111000: out_v[293] = 10'b0111011100;
    16'b0000100100001000: out_v[293] = 10'b0011101011;
    16'b0100000100011000: out_v[293] = 10'b0001011100;
    16'b0001100100010000: out_v[293] = 10'b0111001100;
    16'b0001101100010000: out_v[293] = 10'b0101110111;
    16'b0001100100111001: out_v[293] = 10'b0000111110;
    16'b1000100010011000: out_v[293] = 10'b1000010101;
    16'b0001100100000000: out_v[293] = 10'b0111110011;
    16'b0100000100011001: out_v[293] = 10'b0011110010;
    16'b0000100000001000: out_v[293] = 10'b1110000010;
    16'b0100100100011001: out_v[293] = 10'b0001111110;
    16'b0001101100011000: out_v[293] = 10'b0111011111;
    16'b0100100100001001: out_v[293] = 10'b0011110010;
    16'b0001100000110000: out_v[293] = 10'b0111100011;
    16'b0001101100000000: out_v[293] = 10'b1001011110;
    16'b0000100010010000: out_v[293] = 10'b1101100001;
    16'b0000100000100000: out_v[293] = 10'b0111101010;
    16'b0000100000011001: out_v[293] = 10'b0110001101;
    16'b0001100100001000: out_v[293] = 10'b0111011110;
    16'b0001101000110000: out_v[293] = 10'b0100011011;
    16'b0000100100011001: out_v[293] = 10'b1110001110;
    16'b0000100000101000: out_v[293] = 10'b1101101110;
    16'b0001101100111000: out_v[293] = 10'b0011101111;
    16'b0000100010100000: out_v[293] = 10'b0111010100;
    16'b1101001010111000: out_v[293] = 10'b1110011111;
    16'b0000000110010000: out_v[293] = 10'b1101101000;
    16'b1000000010100000: out_v[293] = 10'b0010101001;
    16'b1001101110111000: out_v[293] = 10'b1000100110;
    16'b0000000000000000: out_v[293] = 10'b1000101000;
    16'b1001100110111000: out_v[293] = 10'b1100101010;
    16'b1101101110111000: out_v[293] = 10'b1001100000;
    16'b0000100110010000: out_v[293] = 10'b1011001111;
    16'b0101000000100000: out_v[293] = 10'b1101100111;
    16'b0000000010000000: out_v[293] = 10'b0010001110;
    16'b1100101110011000: out_v[293] = 10'b1011100110;
    16'b0100101100001000: out_v[293] = 10'b0110111010;
    16'b0000001100010000: out_v[293] = 10'b0011000111;
    16'b0100001110010000: out_v[293] = 10'b1001010001;
    16'b0000101100010000: out_v[293] = 10'b0111001011;
    16'b1100001110011000: out_v[293] = 10'b1111000101;
    16'b0100101100011000: out_v[293] = 10'b0110110111;
    16'b0100001000010000: out_v[293] = 10'b0110110010;
    16'b0000101100001000: out_v[293] = 10'b0011111010;
    16'b0100001100011000: out_v[293] = 10'b1101001110;
    16'b0000001100011000: out_v[293] = 10'b1011000000;
    16'b1000000110011000: out_v[293] = 10'b1001000111;
    16'b0000001110010000: out_v[293] = 10'b0111010001;
    16'b0000101110010000: out_v[293] = 10'b1100101101;
    16'b0000001100000000: out_v[293] = 10'b1100010101;
    16'b0110000100011000: out_v[293] = 10'b1011011010;
    16'b0000101110000000: out_v[293] = 10'b1101011110;
    16'b1000001110011000: out_v[293] = 10'b1001101101;
    16'b0001100110101001: out_v[293] = 10'b0111010001;
    16'b1001101110000000: out_v[293] = 10'b1011011010;
    16'b1001100110100000: out_v[293] = 10'b1101010111;
    16'b1000100010100000: out_v[293] = 10'b1100110101;
    16'b1001101110100000: out_v[293] = 10'b0010100101;
    16'b0001100110000000: out_v[293] = 10'b0111101011;
    16'b1000101110100000: out_v[293] = 10'b1001010001;
    16'b0000100010000000: out_v[293] = 10'b0100111101;
    16'b0000101010100000: out_v[293] = 10'b0011110010;
    16'b1000100010101000: out_v[293] = 10'b1011110101;
    16'b1000101010110000: out_v[293] = 10'b1011000010;
    16'b1000100010001000: out_v[293] = 10'b0111101011;
    16'b1001101010100000: out_v[293] = 10'b0101000100;
    16'b1000101010100000: out_v[293] = 10'b1111100100;
    16'b0001100110100000: out_v[293] = 10'b0101010111;
    16'b1000001010010000: out_v[293] = 10'b0011000101;
    16'b0000000110100000: out_v[293] = 10'b0010110110;
    16'b0001000110000000: out_v[293] = 10'b1111011100;
    16'b0000000110000000: out_v[293] = 10'b0111011001;
    16'b0000100010101000: out_v[293] = 10'b1101001111;
    16'b0001000110100000: out_v[293] = 10'b1001011111;
    16'b0000100110100000: out_v[293] = 10'b0001111110;
    16'b1001101010110000: out_v[293] = 10'b1101001111;
    16'b1001100110000000: out_v[293] = 10'b1100011010;
    16'b1000101010101000: out_v[293] = 10'b1011001010;
    16'b1001000110110000: out_v[293] = 10'b0111110000;
    16'b0000001000110000: out_v[293] = 10'b0100011111;
    16'b0101100100110000: out_v[293] = 10'b0110100011;
    16'b1000001000110000: out_v[293] = 10'b0011101001;
    16'b0001001000110000: out_v[293] = 10'b1110001101;
    16'b0001101100110000: out_v[293] = 10'b0110000100;
    16'b1001001000110000: out_v[293] = 10'b0110001100;
    16'b0001001100110000: out_v[293] = 10'b1110001011;
    16'b0101001000110000: out_v[293] = 10'b0111011000;
    16'b0101101100110000: out_v[293] = 10'b1010101011;
    16'b1101101010111000: out_v[293] = 10'b0101011110;
    16'b0001100100110000: out_v[293] = 10'b1111001000;
    16'b1000101110111000: out_v[293] = 10'b1011001011;
    16'b1000100010111000: out_v[293] = 10'b1101001011;
    16'b1001100110011000: out_v[293] = 10'b0110001011;
    16'b1001101110011000: out_v[293] = 10'b1011100111;
    16'b1100101110011001: out_v[293] = 10'b1111000110;
    16'b1000100110111000: out_v[293] = 10'b0101001010;
    16'b1100101110001000: out_v[293] = 10'b1100000101;
    16'b1000101110001000: out_v[293] = 10'b1100101111;
    16'b1000101010111000: out_v[293] = 10'b1010000111;
    16'b1000101110011000: out_v[293] = 10'b1111110110;
    16'b1100001110011001: out_v[293] = 10'b0110010111;
    16'b1100101110001001: out_v[293] = 10'b1101101010;
    16'b1001101110001000: out_v[293] = 10'b0111100110;
    16'b1001100110010000: out_v[293] = 10'b1111000100;
    default: out_v[293] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100000010000000: out_v[294] = 10'b1101100011;
    16'b0100000110000000: out_v[294] = 10'b1000110000;
    16'b0100100110010100: out_v[294] = 10'b1000010000;
    16'b0100000110000001: out_v[294] = 10'b1000000101;
    16'b0001100010010100: out_v[294] = 10'b0011011101;
    16'b0100100100000100: out_v[294] = 10'b1011011001;
    16'b0001000010010000: out_v[294] = 10'b0001001111;
    16'b0100000010000001: out_v[294] = 10'b0001011001;
    16'b0100100110000000: out_v[294] = 10'b1010011100;
    16'b0100100010000000: out_v[294] = 10'b0001110000;
    16'b0100000010010100: out_v[294] = 10'b1101100101;
    16'b0100000010010000: out_v[294] = 10'b0000111011;
    16'b0100100110000100: out_v[294] = 10'b1001011010;
    16'b0100000100000000: out_v[294] = 10'b1011110001;
    16'b0100100010000100: out_v[294] = 10'b1110110000;
    16'b0100100100000000: out_v[294] = 10'b0100011011;
    16'b0101100110010100: out_v[294] = 10'b1011000001;
    16'b0100000100000001: out_v[294] = 10'b1011010100;
    16'b0001100010000100: out_v[294] = 10'b1011011011;
    16'b0000100010000100: out_v[294] = 10'b1111000010;
    16'b0000000010000000: out_v[294] = 10'b1101001101;
    16'b0001100000010100: out_v[294] = 10'b0000110011;
    16'b0100100010010100: out_v[294] = 10'b1100000000;
    16'b0001000010000000: out_v[294] = 10'b0000010100;
    16'b0100100010010101: out_v[294] = 10'b0101111100;
    16'b0100000000000000: out_v[294] = 10'b0110010111;
    16'b0100100010000101: out_v[294] = 10'b1011111100;
    16'b0100100110000001: out_v[294] = 10'b1111011110;
    16'b0100100110010101: out_v[294] = 10'b0010111011;
    16'b0000000010000001: out_v[294] = 10'b1011010111;
    16'b0001000010010100: out_v[294] = 10'b0000111100;
    16'b0101100010010100: out_v[294] = 10'b1010100011;
    16'b0001100010010101: out_v[294] = 10'b1000011011;
    16'b0100100110000101: out_v[294] = 10'b0110000111;
    16'b0100100010000001: out_v[294] = 10'b1000011110;
    16'b0000000010010000: out_v[294] = 10'b0101001001;
    16'b0000000100000001: out_v[294] = 10'b1111101001;
    16'b0100000110010000: out_v[294] = 10'b1001110111;
    16'b0001000000010000: out_v[294] = 10'b1001011010;
    16'b0000100010010100: out_v[294] = 10'b0011011011;
    16'b0000000100000000: out_v[294] = 10'b1100100101;
    16'b0100000110010100: out_v[294] = 10'b1011100100;
    16'b0100100100000001: out_v[294] = 10'b0000101111;
    16'b0001000000010100: out_v[294] = 10'b0110101011;
    16'b0000000000000001: out_v[294] = 10'b1100000011;
    16'b0000000000000000: out_v[294] = 10'b1100100010;
    16'b0000000100010000: out_v[294] = 10'b0110011011;
    16'b0000000000010000: out_v[294] = 10'b1000110100;
    16'b0001000110000000: out_v[294] = 10'b0010010011;
    16'b0001000110010000: out_v[294] = 10'b1010100110;
    16'b0000000110000001: out_v[294] = 10'b0001010111;
    16'b0001000010010001: out_v[294] = 10'b1010111100;
    16'b0101000110000000: out_v[294] = 10'b1100100100;
    16'b0000000110010000: out_v[294] = 10'b1110100000;
    16'b0001000110000001: out_v[294] = 10'b1001101111;
    16'b0101000100010000: out_v[294] = 10'b1100100101;
    16'b0100000100010000: out_v[294] = 10'b0011000111;
    16'b0100000110010001: out_v[294] = 10'b1111011010;
    16'b0000000110010001: out_v[294] = 10'b1111011011;
    16'b0000000110000000: out_v[294] = 10'b0010111010;
    16'b0101100110010000: out_v[294] = 10'b0111100110;
    16'b0101000000010000: out_v[294] = 10'b0101111010;
    16'b0101000110010000: out_v[294] = 10'b0000010101;
    16'b0001000110010001: out_v[294] = 10'b0011100111;
    16'b0101000110010001: out_v[294] = 10'b0010111111;
    16'b0000000000010001: out_v[294] = 10'b1011010101;
    16'b0101000110000001: out_v[294] = 10'b1011001010;
    16'b0100000000010000: out_v[294] = 10'b0111000110;
    16'b0000000010010001: out_v[294] = 10'b1101110001;
    16'b0001000010000001: out_v[294] = 10'b0010110101;
    16'b0100000100010001: out_v[294] = 10'b1010010100;
    16'b0101000010010000: out_v[294] = 10'b0101001000;
    16'b0100000010110000: out_v[294] = 10'b1100000110;
    16'b0100000010010001: out_v[294] = 10'b0010110000;
    16'b0101000010000000: out_v[294] = 10'b1001000011;
    16'b0000000100100000: out_v[294] = 10'b0011111110;
    16'b0100000110110000: out_v[294] = 10'b1110100011;
    16'b0100000000000001: out_v[294] = 10'b1000011101;
    16'b0000000100000100: out_v[294] = 10'b0101001001;
    16'b0000000100010100: out_v[294] = 10'b1100010010;
    16'b0100000100000100: out_v[294] = 10'b0010010100;
    16'b0100100100010100: out_v[294] = 10'b1011111010;
    16'b0100100000000000: out_v[294] = 10'b1110001111;
    16'b0100000010000100: out_v[294] = 10'b0101011101;
    16'b0000100100000000: out_v[294] = 10'b1111001001;
    16'b0100000100010100: out_v[294] = 10'b1000010111;
    16'b0000100100000100: out_v[294] = 10'b1001100111;
    16'b0000100000000000: out_v[294] = 10'b1100100010;
    16'b0101000010010001: out_v[294] = 10'b0110110111;
    16'b0101000000010100: out_v[294] = 10'b1110100001;
    16'b0101000010010100: out_v[294] = 10'b0100110110;
    16'b0000000100001000: out_v[294] = 10'b1011110101;
    16'b0000001100000000: out_v[294] = 10'b0000100101;
    16'b0101000110010100: out_v[294] = 10'b0111101100;
    16'b0101000010000001: out_v[294] = 10'b1111001001;
    16'b0001100110010100: out_v[294] = 10'b0111011011;
    16'b0001000110010100: out_v[294] = 10'b0000111101;
    16'b0100000110000100: out_v[294] = 10'b0010101111;
    16'b0000000000000100: out_v[294] = 10'b1110001110;
    16'b0000000110010100: out_v[294] = 10'b0111001011;
    default: out_v[294] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000110011000000: out_v[295] = 10'b0110001101;
    16'b0100110011000000: out_v[295] = 10'b1000000101;
    16'b0100100011000000: out_v[295] = 10'b1101110000;
    16'b0100100001000000: out_v[295] = 10'b1000000011;
    16'b0000100011000000: out_v[295] = 10'b0101010100;
    16'b0100000010000000: out_v[295] = 10'b0100011011;
    16'b0100000011000000: out_v[295] = 10'b1110101001;
    16'b0100000001000000: out_v[295] = 10'b0110010101;
    16'b0000010011000000: out_v[295] = 10'b1000100001;
    16'b0100001011000000: out_v[295] = 10'b0000111000;
    16'b0100111011000000: out_v[295] = 10'b1111001111;
    16'b0000100000000000: out_v[295] = 10'b1111100110;
    16'b0100010011000000: out_v[295] = 10'b1001001001;
    16'b0100110001000000: out_v[295] = 10'b1010010101;
    16'b0100100010000000: out_v[295] = 10'b0001000111;
    16'b0000110001000000: out_v[295] = 10'b1010110010;
    16'b0000100001000000: out_v[295] = 10'b0100001001;
    16'b0100101011000000: out_v[295] = 10'b0100000001;
    16'b0000000011000000: out_v[295] = 10'b0010101111;
    16'b0100000000000000: out_v[295] = 10'b1000001101;
    16'b0100010010000000: out_v[295] = 10'b0101110011;
    16'b0000110010000000: out_v[295] = 10'b1010011010;
    16'b0100011011000000: out_v[295] = 10'b0110101000;
    16'b0000111011000000: out_v[295] = 10'b1111000000;
    16'b0000000001000000: out_v[295] = 10'b0001100101;
    16'b0000100010000000: out_v[295] = 10'b0110011000;
    16'b0100110010000000: out_v[295] = 10'b1000111010;
    16'b0000010001000000: out_v[295] = 10'b1111110001;
    16'b0000011011000000: out_v[295] = 10'b0111111011;
    16'b0100100000000000: out_v[295] = 10'b1010110110;
    16'b0000001001000000: out_v[295] = 10'b1100100110;
    16'b0000001000000000: out_v[295] = 10'b1000111010;
    16'b0000000000000000: out_v[295] = 10'b0111101010;
    16'b0000000010000000: out_v[295] = 10'b0111101010;
    16'b0000001010000000: out_v[295] = 10'b0111010100;
    16'b0000001011000000: out_v[295] = 10'b1111000011;
    16'b0100010001000000: out_v[295] = 10'b0011000110;
    16'b0000011000000000: out_v[295] = 10'b1010010011;
    16'b0100001001000000: out_v[295] = 10'b0101011100;
    16'b0000011001000000: out_v[295] = 10'b0111001010;
    16'b0100111001000000: out_v[295] = 10'b0111010110;
    16'b0100010000000000: out_v[295] = 10'b1101111111;
    16'b0100011001000000: out_v[295] = 10'b1010101000;
    16'b0000101001000000: out_v[295] = 10'b1101001101;
    16'b0100110000000000: out_v[295] = 10'b0010011111;
    16'b0100001000000000: out_v[295] = 10'b0110100100;
    16'b0100001010000000: out_v[295] = 10'b0000111110;
    16'b0100011000000000: out_v[295] = 10'b1000001100;
    16'b0100101000000000: out_v[295] = 10'b1101110001;
    16'b0100011010000000: out_v[295] = 10'b0000110010;
    16'b0000010000000000: out_v[295] = 10'b1100110000;
    16'b0000010010000000: out_v[295] = 10'b0110111010;
    16'b0100101001000000: out_v[295] = 10'b1101010010;
    16'b0100111000000000: out_v[295] = 10'b1110010111;
    16'b0000011010000000: out_v[295] = 10'b0100011011;
    16'b0000001011001000: out_v[295] = 10'b1111001001;
    16'b0000001001001000: out_v[295] = 10'b0011100011;
    16'b0000111001000000: out_v[295] = 10'b0101011011;
    16'b0000011001001000: out_v[295] = 10'b0110001011;
    16'b0000101011000000: out_v[295] = 10'b1110101001;
    16'b0000011000001000: out_v[295] = 10'b0101111011;
    16'b0000111000000000: out_v[295] = 10'b0001011101;
    16'b0000110000001000: out_v[295] = 10'b0100111000;
    16'b0000110000000000: out_v[295] = 10'b0010011010;
    16'b0000111010000000: out_v[295] = 10'b1100100011;
    16'b0000101000000000: out_v[295] = 10'b1001111010;
    16'b0000011010101000: out_v[295] = 10'b0111110011;
    16'b0000111010001000: out_v[295] = 10'b1011101100;
    16'b0000011010001000: out_v[295] = 10'b0011101001;
    16'b0000010010001000: out_v[295] = 10'b1100001100;
    16'b0000001010001000: out_v[295] = 10'b1010001111;
    16'b0000110010001000: out_v[295] = 10'b0110110010;
    16'b0000110011001000: out_v[295] = 10'b0111110110;
    16'b0000110001001000: out_v[295] = 10'b0110110100;
    16'b0000111011001000: out_v[295] = 10'b1010111010;
    16'b0000110010101000: out_v[295] = 10'b0001011111;
    16'b0000101010000000: out_v[295] = 10'b1011010010;
    16'b0100101010000000: out_v[295] = 10'b1100010001;
    16'b0000001000100000: out_v[295] = 10'b1001100001;
    16'b0000001010100000: out_v[295] = 10'b1111000100;
    16'b0000011000100000: out_v[295] = 10'b1100100111;
    16'b0000011010100000: out_v[295] = 10'b0111110010;
    default: out_v[295] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000001000101: out_v[296] = 10'b1001100011;
    16'b0000010010000100: out_v[296] = 10'b1101000001;
    16'b1010010011000100: out_v[296] = 10'b0001101010;
    16'b0010010011000100: out_v[296] = 10'b0001100011;
    16'b0000010011000100: out_v[296] = 10'b1001001001;
    16'b0000010010000001: out_v[296] = 10'b1010001111;
    16'b0000010011000000: out_v[296] = 10'b1100110101;
    16'b1010010011000000: out_v[296] = 10'b0110001011;
    16'b0000010010010100: out_v[296] = 10'b0100001111;
    16'b0000010010010000: out_v[296] = 10'b0110100100;
    16'b0000010010010101: out_v[296] = 10'b0011001101;
    16'b0000010010000000: out_v[296] = 10'b1001001101;
    16'b0000010001000100: out_v[296] = 10'b0010011111;
    16'b0000010011000101: out_v[296] = 10'b0101011011;
    16'b0000000001000100: out_v[296] = 10'b0011100000;
    16'b0010010011000101: out_v[296] = 10'b1110000100;
    16'b0000010011010101: out_v[296] = 10'b1110000110;
    16'b0010010011000000: out_v[296] = 10'b0110011101;
    16'b0000010000000100: out_v[296] = 10'b1010011011;
    16'b0000000011000000: out_v[296] = 10'b1001100010;
    16'b1010000001000101: out_v[296] = 10'b1000110101;
    16'b1010010011000101: out_v[296] = 10'b1000001111;
    16'b0000010011010100: out_v[296] = 10'b0111011110;
    16'b1010010001000101: out_v[296] = 10'b0011010110;
    16'b0000000000000000: out_v[296] = 10'b0011011011;
    16'b0010000001000101: out_v[296] = 10'b1111001111;
    16'b0000000000000100: out_v[296] = 10'b1010000000;
    16'b0000000010000100: out_v[296] = 10'b0001110101;
    16'b0000000000010101: out_v[296] = 10'b0001010111;
    16'b0010010001000101: out_v[296] = 10'b1000110110;
    16'b0000000010000000: out_v[296] = 10'b1000011000;
    16'b0010000001000100: out_v[296] = 10'b1010100111;
    16'b0010010001000100: out_v[296] = 10'b1101000110;
    16'b0000000011000100: out_v[296] = 10'b1101111000;
    16'b0000010010000101: out_v[296] = 10'b0001100110;
    16'b0000000001010101: out_v[296] = 10'b0011011111;
    16'b0010000001010101: out_v[296] = 10'b0111011000;
    16'b0000000000010001: out_v[296] = 10'b0001000011;
    16'b0000000001000000: out_v[296] = 10'b0111110111;
    16'b0000000000010000: out_v[296] = 10'b1100110100;
    16'b0000000000000001: out_v[296] = 10'b1111011001;
    16'b0000000010010001: out_v[296] = 10'b0000110100;
    16'b0000000001010000: out_v[296] = 10'b1001111010;
    16'b0010000001000000: out_v[296] = 10'b1011001011;
    16'b0010000001010000: out_v[296] = 10'b1000101111;
    16'b0000000010000001: out_v[296] = 10'b1100011010;
    16'b0000010010010001: out_v[296] = 10'b1011000010;
    16'b0000000001010001: out_v[296] = 10'b0111010001;
    16'b1010000001000001: out_v[296] = 10'b1110101100;
    16'b1010000000010001: out_v[296] = 10'b0100110011;
    16'b0010010011010100: out_v[296] = 10'b1110010110;
    16'b0010000001000001: out_v[296] = 10'b0000110101;
    16'b1010000011010001: out_v[296] = 10'b1001111001;
    16'b1010000001000000: out_v[296] = 10'b1010000100;
    16'b1010010010010001: out_v[296] = 10'b0011110110;
    16'b0010000001010001: out_v[296] = 10'b0111010000;
    16'b1010000000000001: out_v[296] = 10'b0100010011;
    16'b0000010011010001: out_v[296] = 10'b0010100111;
    16'b1010010010000001: out_v[296] = 10'b1111011100;
    16'b0000010000010001: out_v[296] = 10'b1010100010;
    16'b0010010011010001: out_v[296] = 10'b1010110101;
    16'b0010000011000101: out_v[296] = 10'b1101110110;
    16'b0000000001000001: out_v[296] = 10'b1001110101;
    16'b1010010011010001: out_v[296] = 10'b1100110001;
    16'b1010010011010101: out_v[296] = 10'b1101011100;
    16'b1010010011010100: out_v[296] = 10'b0101010110;
    16'b0000010011000001: out_v[296] = 10'b1001110000;
    16'b1010010010000101: out_v[296] = 10'b0011001110;
    16'b1010000010000001: out_v[296] = 10'b1010111001;
    16'b0000000011000101: out_v[296] = 10'b1010000100;
    16'b0000000011000001: out_v[296] = 10'b0010110100;
    16'b1010000011000001: out_v[296] = 10'b1010110110;
    16'b1010000001010001: out_v[296] = 10'b1110000101;
    16'b0010010011000001: out_v[296] = 10'b0011111011;
    16'b0000000010000101: out_v[296] = 10'b0100000110;
    16'b0010010011010101: out_v[296] = 10'b0101010010;
    16'b0000000010010101: out_v[296] = 10'b0010000100;
    16'b1010010011000001: out_v[296] = 10'b0111110011;
    16'b0010000011000001: out_v[296] = 10'b1011011111;
    16'b1010000011000101: out_v[296] = 10'b1010010110;
    16'b0010000011010001: out_v[296] = 10'b1111010001;
    16'b1010010001010001: out_v[296] = 10'b1011101010;
    16'b0010010011010000: out_v[296] = 10'b1100000101;
    16'b0000000010010000: out_v[296] = 10'b0010101000;
    16'b1010000011010000: out_v[296] = 10'b1010010101;
    16'b1010000001010000: out_v[296] = 10'b1001101010;
    16'b1010000011000100: out_v[296] = 10'b1001100110;
    16'b1010000000010000: out_v[296] = 10'b1100001011;
    16'b0010000011010000: out_v[296] = 10'b0000111111;
    16'b1010000000000000: out_v[296] = 10'b1101100100;
    16'b0000000001011000: out_v[296] = 10'b1000101011;
    16'b0000010011010000: out_v[296] = 10'b1000111011;
    16'b1010000011010100: out_v[296] = 10'b0011111001;
    16'b1010000001010100: out_v[296] = 10'b0100100000;
    16'b0000000001010100: out_v[296] = 10'b1000110010;
    16'b0000000010010100: out_v[296] = 10'b0010101011;
    16'b1010010011010000: out_v[296] = 10'b1101010101;
    16'b0010000001011000: out_v[296] = 10'b0001110111;
    16'b0000000011010100: out_v[296] = 10'b1000001110;
    16'b1010000010000000: out_v[296] = 10'b1111110011;
    16'b0010000011000000: out_v[296] = 10'b0001001011;
    16'b1010000001011000: out_v[296] = 10'b0001011111;
    16'b1010000010010000: out_v[296] = 10'b0110110111;
    16'b0010000000010000: out_v[296] = 10'b1111001001;
    16'b0010000000000000: out_v[296] = 10'b0011001110;
    16'b0000000011010000: out_v[296] = 10'b0000011001;
    16'b0010000011010100: out_v[296] = 10'b1010111100;
    16'b1010000011000000: out_v[296] = 10'b1011110011;
    16'b0010000001010100: out_v[296] = 10'b0100011010;
    16'b0000000001011100: out_v[296] = 10'b1000010011;
    16'b0000000000010100: out_v[296] = 10'b1000010010;
    16'b0000010000000101: out_v[296] = 10'b1000101010;
    16'b1000000000010100: out_v[296] = 10'b0000011101;
    16'b1010000000010100: out_v[296] = 10'b0001111011;
    16'b0000010000000001: out_v[296] = 10'b0000111010;
    16'b0000010001000101: out_v[296] = 10'b1000010011;
    16'b1000000000010000: out_v[296] = 10'b0100011011;
    16'b1000000000000001: out_v[296] = 10'b0001111111;
    16'b0000010001000001: out_v[296] = 10'b0110110010;
    16'b0000010000010100: out_v[296] = 10'b1001110110;
    16'b0000010000010000: out_v[296] = 10'b0001101110;
    16'b0000000000000101: out_v[296] = 10'b0110001010;
    16'b0000010000000000: out_v[296] = 10'b1111001000;
    16'b1010000000010101: out_v[296] = 10'b0111000010;
    16'b0000010001010001: out_v[296] = 10'b1111101110;
    16'b1010000000000101: out_v[296] = 10'b0100111010;
    16'b0000010001010101: out_v[296] = 10'b1001001110;
    16'b1000000000000101: out_v[296] = 10'b0011101011;
    16'b0010010001010101: out_v[296] = 10'b1011111011;
    16'b0000010000010101: out_v[296] = 10'b0111100100;
    16'b1010000001010101: out_v[296] = 10'b1100000100;
    16'b0000000000001100: out_v[296] = 10'b0011001101;
    16'b0000000001001000: out_v[296] = 10'b0111101101;
    16'b0000000000001000: out_v[296] = 10'b0111000010;
    16'b1010000001000100: out_v[296] = 10'b1010110111;
    16'b1010000001001100: out_v[296] = 10'b0110101011;
    16'b0000000001001100: out_v[296] = 10'b0011110111;
    16'b1010000001001000: out_v[296] = 10'b1111110011;
    16'b0010000001001000: out_v[296] = 10'b0011110101;
    16'b0000000011010101: out_v[296] = 10'b1110011010;
    16'b0000000001011101: out_v[296] = 10'b0111011011;
    16'b0000000011010001: out_v[296] = 10'b1100101100;
    16'b0010000011010101: out_v[296] = 10'b1110011011;
    16'b0000000000001101: out_v[296] = 10'b1100001100;
    16'b0000000000011100: out_v[296] = 10'b1100101010;
    16'b0000000000011000: out_v[296] = 10'b1011100101;
    16'b0000000001001101: out_v[296] = 10'b1101011010;
    default: out_v[296] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0011110000010010: out_v[297] = 10'b0010001001;
    16'b0000110010000010: out_v[297] = 10'b1010011101;
    16'b1010110010000010: out_v[297] = 10'b1111010110;
    16'b1011110010000010: out_v[297] = 10'b0000110110;
    16'b0000110000010010: out_v[297] = 10'b1001000110;
    16'b1010110000000000: out_v[297] = 10'b0110010001;
    16'b1011110010000000: out_v[297] = 10'b0001110001;
    16'b0011110000000010: out_v[297] = 10'b1010100111;
    16'b0000110010010010: out_v[297] = 10'b1101011110;
    16'b1000110010000010: out_v[297] = 10'b1110100011;
    16'b0000111010010010: out_v[297] = 10'b0011010001;
    16'b0011110010010010: out_v[297] = 10'b0011101000;
    16'b0010110010000010: out_v[297] = 10'b1111100101;
    16'b0001110010000010: out_v[297] = 10'b0000011110;
    16'b0001110000010010: out_v[297] = 10'b1101000111;
    16'b0011110010000010: out_v[297] = 10'b1010110110;
    16'b1000110000000010: out_v[297] = 10'b1100010011;
    16'b1010110010000000: out_v[297] = 10'b1101001001;
    16'b0000001010000010: out_v[297] = 10'b0001001101;
    16'b0011110010000000: out_v[297] = 10'b1011011011;
    16'b0000110000000010: out_v[297] = 10'b1110110000;
    16'b0001110010010010: out_v[297] = 10'b1010111011;
    16'b0011000000010010: out_v[297] = 10'b1111000011;
    16'b0011100000010010: out_v[297] = 10'b0001000011;
    16'b1011111010010010: out_v[297] = 10'b0111100111;
    16'b1000001010000010: out_v[297] = 10'b0111000001;
    16'b0010110000010010: out_v[297] = 10'b0111010011;
    16'b1010110000010000: out_v[297] = 10'b1000101111;
    16'b1011100010000000: out_v[297] = 10'b0001110111;
    16'b1000111010000010: out_v[297] = 10'b1111001110;
    16'b1010111010000010: out_v[297] = 10'b1001111111;
    16'b1011110010010010: out_v[297] = 10'b0111110000;
    16'b0001110000010000: out_v[297] = 10'b1100100101;
    16'b0000001010010010: out_v[297] = 10'b1011001111;
    16'b1010111010010010: out_v[297] = 10'b0011001111;
    16'b1001110010000000: out_v[297] = 10'b0010101011;
    16'b0011111010010010: out_v[297] = 10'b1010111011;
    16'b0010110010010010: out_v[297] = 10'b0100110111;
    16'b1000001010010010: out_v[297] = 10'b1010110100;
    16'b0000001010010000: out_v[297] = 10'b0101010001;
    16'b0000001000000000: out_v[297] = 10'b1001010110;
    16'b0001001000000000: out_v[297] = 10'b0111100011;
    16'b0001101000000000: out_v[297] = 10'b1011100111;
    16'b0000101000000000: out_v[297] = 10'b1010000110;
    16'b0000000000000000: out_v[297] = 10'b0010111001;
    16'b0000000000010000: out_v[297] = 10'b0001001011;
    16'b0001111000000000: out_v[297] = 10'b1001100111;
    16'b0000000010010000: out_v[297] = 10'b1000101010;
    16'b0000111000000000: out_v[297] = 10'b0101110111;
    16'b0000001000010000: out_v[297] = 10'b0000111011;
    16'b0001111000010000: out_v[297] = 10'b0110011100;
    16'b0001111010010000: out_v[297] = 10'b0001111110;
    16'b0001111010000010: out_v[297] = 10'b1010101111;
    16'b0001001010010000: out_v[297] = 10'b0111011100;
    16'b0001011010010000: out_v[297] = 10'b1000010000;
    16'b0001110010010000: out_v[297] = 10'b1101010000;
    16'b0001001010000000: out_v[297] = 10'b1101111000;
    16'b1000001000010010: out_v[297] = 10'b0111010010;
    16'b0001100010010000: out_v[297] = 10'b1000110101;
    16'b0001001000010000: out_v[297] = 10'b1100000011;
    16'b0001000000010000: out_v[297] = 10'b1010010111;
    16'b0001110000000000: out_v[297] = 10'b1100011101;
    16'b0001100000010000: out_v[297] = 10'b0001011101;
    16'b0000111010010000: out_v[297] = 10'b1000110110;
    16'b1001111000010000: out_v[297] = 10'b0110100011;
    16'b0011111010010000: out_v[297] = 10'b1000011110;
    16'b0001111010000000: out_v[297] = 10'b1011111011;
    16'b0001011000010000: out_v[297] = 10'b1010011110;
    16'b1001001000010010: out_v[297] = 10'b0011101100;
    16'b0001001010010010: out_v[297] = 10'b1010111011;
    16'b1001111010010000: out_v[297] = 10'b1100011010;
    16'b0011111000010000: out_v[297] = 10'b0100111010;
    16'b0010001000010000: out_v[297] = 10'b1010100101;
    16'b1001001010000010: out_v[297] = 10'b1101110111;
    16'b0001111010010010: out_v[297] = 10'b0010111010;
    16'b1001001010010000: out_v[297] = 10'b0110011111;
    16'b1000000000010010: out_v[297] = 10'b0100101101;
    16'b0000111000010000: out_v[297] = 10'b1011111001;
    16'b1001011010010000: out_v[297] = 10'b0001100011;
    16'b0011001010010000: out_v[297] = 10'b1111000111;
    16'b0001001000010010: out_v[297] = 10'b1110101110;
    16'b0001001010000010: out_v[297] = 10'b1010000101;
    16'b0000011000010000: out_v[297] = 10'b0001011100;
    16'b1001111010010010: out_v[297] = 10'b1010111110;
    16'b0000110000010000: out_v[297] = 10'b0111010101;
    16'b0000110010010000: out_v[297] = 10'b1110110101;
    16'b0001000010010000: out_v[297] = 10'b1000000100;
    16'b0000011010010000: out_v[297] = 10'b1001011100;
    16'b1001001010010010: out_v[297] = 10'b1000100101;
    16'b0001111000010010: out_v[297] = 10'b1000110101;
    16'b0000001000010010: out_v[297] = 10'b1010011001;
    16'b0011011010010000: out_v[297] = 10'b1001001110;
    16'b0001011000010010: out_v[297] = 10'b0101100110;
    16'b0001110000000010: out_v[297] = 10'b0100001110;
    16'b0001110010000000: out_v[297] = 10'b1011001011;
    16'b0001110000000100: out_v[297] = 10'b1110010100;
    16'b0001100000000000: out_v[297] = 10'b1100111100;
    16'b0000110000100000: out_v[297] = 10'b0000100110;
    16'b0000110000100010: out_v[297] = 10'b0110101010;
    16'b0001000000000000: out_v[297] = 10'b0010111101;
    16'b0001110000000110: out_v[297] = 10'b0101011011;
    16'b0001000000000010: out_v[297] = 10'b1101011001;
    16'b0011110000000000: out_v[297] = 10'b1001001111;
    16'b0000110010000000: out_v[297] = 10'b0010001100;
    16'b0001100010000010: out_v[297] = 10'b1100110011;
    16'b0001100010000000: out_v[297] = 10'b0111011001;
    16'b0001100000000010: out_v[297] = 10'b0010111101;
    16'b1001110010000010: out_v[297] = 10'b0101010110;
    16'b0000110000000000: out_v[297] = 10'b1111000000;
    16'b0001000010000000: out_v[297] = 10'b1010011001;
    16'b0010110000000000: out_v[297] = 10'b1001111101;
    16'b0010111000010010: out_v[297] = 10'b1100011000;
    16'b0000001000100010: out_v[297] = 10'b0011000010;
    16'b0010110000000010: out_v[297] = 10'b1101110110;
    16'b0000000000000010: out_v[297] = 10'b1000010001;
    16'b0010001000000010: out_v[297] = 10'b1001011111;
    16'b0010010000000010: out_v[297] = 10'b1110100111;
    16'b0011001000000010: out_v[297] = 10'b1000011111;
    16'b0000001000000010: out_v[297] = 10'b0010000111;
    16'b0000100000000010: out_v[297] = 10'b0100110101;
    16'b0001001000000010: out_v[297] = 10'b0000001011;
    16'b0010111000000010: out_v[297] = 10'b0111011001;
    16'b0010000000000010: out_v[297] = 10'b0000110011;
    16'b0010001000100010: out_v[297] = 10'b1001010010;
    16'b0010100000000010: out_v[297] = 10'b1011100110;
    16'b0000111000010010: out_v[297] = 10'b1001111010;
    16'b1010001000000010: out_v[297] = 10'b1110101101;
    16'b0010001000010010: out_v[297] = 10'b0100011100;
    16'b0010101000010010: out_v[297] = 10'b0100110011;
    16'b0000010000000010: out_v[297] = 10'b0011111011;
    16'b1000001000000010: out_v[297] = 10'b1100101001;
    16'b0011111000010010: out_v[297] = 10'b1011010000;
    16'b1010110000000010: out_v[297] = 10'b0110001000;
    16'b0000101000010010: out_v[297] = 10'b1101011001;
    16'b1010111000010010: out_v[297] = 10'b1010000011;
    16'b0010101000000010: out_v[297] = 10'b0111001101;
    16'b0000111000000010: out_v[297] = 10'b0111000010;
    16'b0000101000000010: out_v[297] = 10'b1100110011;
    16'b0000001010000000: out_v[297] = 10'b0110011100;
    16'b0000000010000010: out_v[297] = 10'b0100111011;
    16'b0010110010000000: out_v[297] = 10'b0000001011;
    16'b1000001000010000: out_v[297] = 10'b0000111010;
    16'b0011000000000010: out_v[297] = 10'b1011100111;
    16'b0010110000100010: out_v[297] = 10'b0000111010;
    16'b0010111010000010: out_v[297] = 10'b1000110111;
    16'b0010111000100010: out_v[297] = 10'b1000000101;
    16'b1000110010000000: out_v[297] = 10'b1001110101;
    16'b0011100000000010: out_v[297] = 10'b1010100010;
    16'b0010011000010010: out_v[297] = 10'b1100110010;
    16'b0011011000010010: out_v[297] = 10'b1011101111;
    16'b0000010000010010: out_v[297] = 10'b1011000011;
    16'b0000011000010010: out_v[297] = 10'b0111111001;
    16'b0000001000100000: out_v[297] = 10'b1011010101;
    16'b0010001000000000: out_v[297] = 10'b0110111001;
    16'b0010001000100000: out_v[297] = 10'b1000101011;
    16'b0010101000100000: out_v[297] = 10'b1101111101;
    16'b0010111000000000: out_v[297] = 10'b0111000100;
    16'b0010110000100000: out_v[297] = 10'b0011111111;
    16'b0010101000000000: out_v[297] = 10'b0111110001;
    16'b0010111000100000: out_v[297] = 10'b0101111110;
    16'b0010010000000000: out_v[297] = 10'b0110111011;
    16'b0010000000100000: out_v[297] = 10'b1111100110;
    16'b0010000000000000: out_v[297] = 10'b0010100100;
    16'b0010101000100010: out_v[297] = 10'b1011100111;
    16'b0010001010010000: out_v[297] = 10'b0011001011;
    16'b0000101000100000: out_v[297] = 10'b1001101001;
    16'b0010001000110000: out_v[297] = 10'b0010101010;
    16'b0000100000000000: out_v[297] = 10'b1110010100;
    16'b0010100000000000: out_v[297] = 10'b0000111000;
    16'b0010100000100000: out_v[297] = 10'b1001000110;
    16'b0000111000100000: out_v[297] = 10'b0001011010;
    16'b0000001000110000: out_v[297] = 10'b1011001001;
    16'b0000000000100000: out_v[297] = 10'b0001101111;
    16'b0010110010010000: out_v[297] = 10'b0001100111;
    16'b0010001010010010: out_v[297] = 10'b0100011010;
    16'b0011110000010000: out_v[297] = 10'b1110110110;
    16'b0011111000000010: out_v[297] = 10'b0110001100;
    16'b0011111000000000: out_v[297] = 10'b0101010111;
    16'b0011110010010000: out_v[297] = 10'b1110010110;
    16'b0010111010010000: out_v[297] = 10'b1010101100;
    16'b0000101010010000: out_v[297] = 10'b1100010110;
    16'b0000101000010000: out_v[297] = 10'b0111111110;
    16'b0011000000010000: out_v[297] = 10'b0100010010;
    16'b0010110000010000: out_v[297] = 10'b1110111010;
    16'b0010111010010010: out_v[297] = 10'b1011110010;
    16'b0001101000010000: out_v[297] = 10'b0101101000;
    16'b0001101010010000: out_v[297] = 10'b0001001010;
    16'b0011100000010000: out_v[297] = 10'b0000111011;
    16'b0000000000100010: out_v[297] = 10'b1010001110;
    16'b0010100000100010: out_v[297] = 10'b1100100111;
    16'b0000001000110010: out_v[297] = 10'b1001101110;
    16'b0010111000010000: out_v[297] = 10'b0001111101;
    16'b0000101000100010: out_v[297] = 10'b0111111011;
    default: out_v[297] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000100100001000: out_v[298] = 10'b0001011011;
    16'b0000000100001000: out_v[298] = 10'b1010000011;
    16'b0010100100001000: out_v[298] = 10'b0010110101;
    16'b0010010100000000: out_v[298] = 10'b0010111101;
    16'b0000000100011000: out_v[298] = 10'b1100110010;
    16'b0000100100001011: out_v[298] = 10'b0101000011;
    16'b0000100110011001: out_v[298] = 10'b1100011001;
    16'b0000010110001000: out_v[298] = 10'b0000011001;
    16'b0010000100001000: out_v[298] = 10'b1000110111;
    16'b0000100100001001: out_v[298] = 10'b1001011110;
    16'b0010010100001000: out_v[298] = 10'b0111000110;
    16'b0000110100001011: out_v[298] = 10'b1110110010;
    16'b0000100000001001: out_v[298] = 10'b0001011011;
    16'b0010100100001001: out_v[298] = 10'b1111101001;
    16'b0010110100001000: out_v[298] = 10'b0011001011;
    16'b0000000100000000: out_v[298] = 10'b1010101001;
    16'b0000110100000000: out_v[298] = 10'b0011010011;
    16'b0010110100001001: out_v[298] = 10'b0001011110;
    16'b0000010100000000: out_v[298] = 10'b1011001111;
    16'b0010110100000000: out_v[298] = 10'b0010001001;
    16'b0000100110001001: out_v[298] = 10'b1110000101;
    16'b0000000110001000: out_v[298] = 10'b1111110010;
    16'b0010100100011001: out_v[298] = 10'b1011100111;
    16'b0000000110011000: out_v[298] = 10'b0000111100;
    16'b0000010100001010: out_v[298] = 10'b0010011011;
    16'b0000110100001000: out_v[298] = 10'b0110001010;
    16'b0000110100001001: out_v[298] = 10'b1000101100;
    16'b0000100010001001: out_v[298] = 10'b0101000110;
    16'b0000010100001000: out_v[298] = 10'b1101101111;
    16'b0000100110001011: out_v[298] = 10'b1110100110;
    16'b0000000100001001: out_v[298] = 10'b1011001110;
    16'b0000000100001010: out_v[298] = 10'b1001011010;
    16'b0000010110000000: out_v[298] = 10'b1001111001;
    16'b0000100100011001: out_v[298] = 10'b0010110001;
    16'b0000010100000010: out_v[298] = 10'b1110100101;
    16'b0010110100000001: out_v[298] = 10'b0011010001;
    16'b0000110100000001: out_v[298] = 10'b0100100101;
    16'b0000110110001011: out_v[298] = 10'b0111101100;
    16'b0000100010011001: out_v[298] = 10'b0011010011;
    16'b0000100100011000: out_v[298] = 10'b1011010111;
    16'b0000100110011011: out_v[298] = 10'b1011001010;
    16'b0000100010000001: out_v[298] = 10'b0010000110;
    16'b0000000110000001: out_v[298] = 10'b0110001000;
    16'b0000000010000001: out_v[298] = 10'b0110110101;
    16'b0010000110000001: out_v[298] = 10'b1110110101;
    16'b0000000110010001: out_v[298] = 10'b1111001100;
    16'b0000100010000000: out_v[298] = 10'b1010101111;
    16'b0010000010000001: out_v[298] = 10'b0111101001;
    16'b0010000110000000: out_v[298] = 10'b0100010010;
    16'b0000100110000001: out_v[298] = 10'b1100110101;
    16'b0010100110000001: out_v[298] = 10'b1000111101;
    16'b0000000010010001: out_v[298] = 10'b1000110011;
    16'b0000000010000000: out_v[298] = 10'b1101100111;
    16'b0000100110010001: out_v[298] = 10'b1101001111;
    16'b0010100110010001: out_v[298] = 10'b1010101011;
    16'b0010000010000000: out_v[298] = 10'b0111100011;
    16'b0000100010010001: out_v[298] = 10'b0001110101;
    16'b0000000110000000: out_v[298] = 10'b1001101010;
    16'b0010000110010001: out_v[298] = 10'b1011011001;
    16'b0000000000000000: out_v[298] = 10'b0010010011;
    16'b0010110110000001: out_v[298] = 10'b1110110011;
    16'b0010101100001001: out_v[298] = 10'b0100111101;
    16'b0010111100000001: out_v[298] = 10'b1101111010;
    16'b0000110110000001: out_v[298] = 10'b1000110100;
    16'b0010000100001001: out_v[298] = 10'b1001001111;
    16'b0010110110011001: out_v[298] = 10'b1011111000;
    16'b0010110100001011: out_v[298] = 10'b1111100001;
    16'b0000100100000001: out_v[298] = 10'b1110100110;
    16'b0010100100000001: out_v[298] = 10'b0011110100;
    16'b0010100110001001: out_v[298] = 10'b1111011000;
    16'b0010111110000001: out_v[298] = 10'b1111010100;
    16'b0010111000000001: out_v[298] = 10'b1011001011;
    16'b0010111100001001: out_v[298] = 10'b0111000110;
    16'b0010101100000001: out_v[298] = 10'b1011111101;
    16'b0000110110010001: out_v[298] = 10'b1010011100;
    16'b0010110110001001: out_v[298] = 10'b0100100111;
    16'b0010111100001011: out_v[298] = 10'b0011111111;
    16'b0000000010001000: out_v[298] = 10'b1010000100;
    16'b0010110110010001: out_v[298] = 10'b0010110100;
    16'b0010010110000000: out_v[298] = 10'b0100011011;
    16'b0010110000000001: out_v[298] = 10'b1111001101;
    16'b0010010100000001: out_v[298] = 10'b1000101111;
    16'b0010110110000000: out_v[298] = 10'b1011011110;
    16'b0010110100011001: out_v[298] = 10'b0011111101;
    16'b0010010100001001: out_v[298] = 10'b0011100100;
    16'b0000110010000001: out_v[298] = 10'b0000110111;
    16'b0010000110011000: out_v[298] = 10'b1101010101;
    16'b0000010100011000: out_v[298] = 10'b1111100110;
    16'b0010110110011000: out_v[298] = 10'b0110010010;
    16'b0010010110011000: out_v[298] = 10'b0111010011;
    16'b0000010110011000: out_v[298] = 10'b1011001100;
    16'b0000000110010000: out_v[298] = 10'b0100011011;
    16'b0000010110010000: out_v[298] = 10'b1001111000;
    16'b0000110110011000: out_v[298] = 10'b1111011110;
    16'b0000010010011000: out_v[298] = 10'b0010011011;
    16'b0010100110011001: out_v[298] = 10'b1111101100;
    16'b0010100110011000: out_v[298] = 10'b1111100110;
    16'b0010000110001000: out_v[298] = 10'b0000111111;
    16'b0000100110011000: out_v[298] = 10'b0111110111;
    16'b0010100110010000: out_v[298] = 10'b0110110100;
    16'b0010000110010000: out_v[298] = 10'b0011001101;
    16'b0010010110010000: out_v[298] = 10'b0100000110;
    16'b0000000110011001: out_v[298] = 10'b1000110110;
    16'b0010110110001000: out_v[298] = 10'b0011011000;
    16'b0000000100010000: out_v[298] = 10'b1011100110;
    16'b0010010110001000: out_v[298] = 10'b0100110011;
    16'b0000110110011001: out_v[298] = 10'b1000001011;
    16'b0000000000001001: out_v[298] = 10'b0111100100;
    16'b0000000010001001: out_v[298] = 10'b0111000011;
    16'b0000000000010001: out_v[298] = 10'b0001010010;
    16'b0000010000001000: out_v[298] = 10'b0010011000;
    16'b0000100000000001: out_v[298] = 10'b1010111011;
    16'b0000000000010000: out_v[298] = 10'b0101111111;
    16'b0000000000001000: out_v[298] = 10'b0110011000;
    16'b0000000000000001: out_v[298] = 10'b1001011010;
    16'b0000000010011000: out_v[298] = 10'b1001111111;
    16'b0000000110001001: out_v[298] = 10'b0010111010;
    16'b0000000000011000: out_v[298] = 10'b0110101110;
    16'b0000000100000001: out_v[298] = 10'b1110101011;
    16'b0000000000001010: out_v[298] = 10'b0111010010;
    16'b0000010000001001: out_v[298] = 10'b0011111010;
    16'b0000010000011000: out_v[298] = 10'b0001111011;
    16'b0000000010010000: out_v[298] = 10'b1001101011;
    16'b0000100000010001: out_v[298] = 10'b1100100100;
    16'b0000000010011001: out_v[298] = 10'b0010011101;
    16'b0000010000001010: out_v[298] = 10'b0111011010;
    16'b0000000000011001: out_v[298] = 10'b0010101011;
    16'b0001100000010001: out_v[298] = 10'b1001111110;
    16'b0001100010010001: out_v[298] = 10'b0010100110;
    16'b0000000100010001: out_v[298] = 10'b1101000001;
    16'b0001000000000001: out_v[298] = 10'b1101001111;
    16'b0001100010000001: out_v[298] = 10'b1110001000;
    16'b0000110100011000: out_v[298] = 10'b0100101000;
    16'b0000010100010000: out_v[298] = 10'b1010001110;
    16'b0001000000000000: out_v[298] = 10'b0101010001;
    16'b0000100100010001: out_v[298] = 10'b0110011011;
    16'b0000100100010000: out_v[298] = 10'b0010011011;
    16'b0010010100011000: out_v[298] = 10'b0110100010;
    16'b0010000100011000: out_v[298] = 10'b1001100111;
    16'b0010110100011000: out_v[298] = 10'b1011010001;
    16'b0000101100001001: out_v[298] = 10'b0110001101;
    16'b0000111100001001: out_v[298] = 10'b0111001110;
    16'b0010100000000001: out_v[298] = 10'b1011101100;
    16'b0000110000001001: out_v[298] = 10'b0111001010;
    16'b0010101100011001: out_v[298] = 10'b1100111011;
    16'b0000101100011001: out_v[298] = 10'b1110000011;
    16'b0000101100010001: out_v[298] = 10'b1011011100;
    16'b0000010000000001: out_v[298] = 10'b1011111011;
    16'b0010000000001001: out_v[298] = 10'b0001001100;
    16'b0000101110011001: out_v[298] = 10'b0011000000;
    16'b0000101100000001: out_v[298] = 10'b0001011000;
    16'b0010100000001001: out_v[298] = 10'b1001101011;
    16'b0000111100011001: out_v[298] = 10'b0111001011;
    16'b0000101010011001: out_v[298] = 10'b1011000110;
    16'b0000101100010000: out_v[298] = 10'b1010011110;
    16'b0000110000000001: out_v[298] = 10'b1101000010;
    16'b0000101100011000: out_v[298] = 10'b1100011101;
    16'b0010101110011001: out_v[298] = 10'b0011011110;
    16'b0010110000001001: out_v[298] = 10'b0010010011;
    16'b0000101110010001: out_v[298] = 10'b0101001101;
    16'b0000101100001000: out_v[298] = 10'b1010111011;
    16'b0010111100011001: out_v[298] = 10'b0110101111;
    16'b0010010000001001: out_v[298] = 10'b0111011010;
    16'b0000101110011000: out_v[298] = 10'b1011100011;
    16'b0010100000011001: out_v[298] = 10'b1110101011;
    16'b0000110010001001: out_v[298] = 10'b0101001101;
    16'b0010100010001001: out_v[298] = 10'b1111100010;
    16'b0010100010011001: out_v[298] = 10'b1111101110;
    16'b0000110010010001: out_v[298] = 10'b1001001000;
    16'b0000100010101001: out_v[298] = 10'b0011011011;
    16'b0000010010001000: out_v[298] = 10'b1001101100;
    16'b0000100000100001: out_v[298] = 10'b0110111011;
    16'b0000100010100001: out_v[298] = 10'b0011111000;
    16'b0000000000100001: out_v[298] = 10'b0110111101;
    16'b0000000000101001: out_v[298] = 10'b1011100110;
    16'b0000000010100001: out_v[298] = 10'b1110101111;
    16'b0000100000101001: out_v[298] = 10'b1000101011;
    16'b0000100110010000: out_v[298] = 10'b0111110000;
    16'b0001000100010001: out_v[298] = 10'b1011001001;
    16'b0010100110000000: out_v[298] = 10'b0101110001;
    16'b0000100110000000: out_v[298] = 10'b0111110011;
    16'b0000100100000000: out_v[298] = 10'b0111010001;
    16'b0010100100010000: out_v[298] = 10'b1011100001;
    16'b0000110110010000: out_v[298] = 10'b0110010001;
    16'b0010000100010000: out_v[298] = 10'b0101011001;
    default: out_v[298] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000100110010000: out_v[299] = 10'b0110111011;
    16'b0000100111010000: out_v[299] = 10'b1010100111;
    16'b0010100111010000: out_v[299] = 10'b0101011101;
    16'b0000000101010001: out_v[299] = 10'b0110111011;
    16'b0000000111010000: out_v[299] = 10'b1011011010;
    16'b0010000011000000: out_v[299] = 10'b0111101100;
    16'b0000100110011000: out_v[299] = 10'b1100000010;
    16'b0000100111011001: out_v[299] = 10'b0010011111;
    16'b0000000111110000: out_v[299] = 10'b1010110000;
    16'b0010000111010000: out_v[299] = 10'b1000111111;
    16'b0000100101011000: out_v[299] = 10'b1001001110;
    16'b0000000101110000: out_v[299] = 10'b1000011111;
    16'b0000100101010001: out_v[299] = 10'b0101110111;
    16'b0000000111000000: out_v[299] = 10'b1000100010;
    16'b0000000110010000: out_v[299] = 10'b0100010001;
    16'b0010100111000000: out_v[299] = 10'b1101100011;
    16'b0010000101000000: out_v[299] = 10'b1110110001;
    16'b0010000111000000: out_v[299] = 10'b0000001001;
    16'b0010100101000000: out_v[299] = 10'b1001101011;
    16'b0010000101010000: out_v[299] = 10'b0010000111;
    16'b0000100101011001: out_v[299] = 10'b0111110111;
    16'b0000000101010000: out_v[299] = 10'b0001011111;
    16'b0010100111010001: out_v[299] = 10'b0111110011;
    16'b0000100111010001: out_v[299] = 10'b1100100011;
    16'b0000000011010000: out_v[299] = 10'b1011101110;
    16'b0000000101110001: out_v[299] = 10'b0010111011;
    16'b0000000101110011: out_v[299] = 10'b1000001111;
    16'b0000000111110010: out_v[299] = 10'b1100001111;
    16'b0000000101000000: out_v[299] = 10'b1000110111;
    16'b0000100100011000: out_v[299] = 10'b1000100011;
    16'b0000000111110001: out_v[299] = 10'b1010111111;
    16'b0000100111011000: out_v[299] = 10'b1100110001;
    16'b0000000111010001: out_v[299] = 10'b1111011000;
    16'b0010000111110000: out_v[299] = 10'b1101011111;
    16'b0000100101010000: out_v[299] = 10'b1101010111;
    16'b0000000100010000: out_v[299] = 10'b1111100101;
    16'b0010000111010001: out_v[299] = 10'b1010000110;
    16'b0000100100011001: out_v[299] = 10'b1011100110;
    16'b0010000111100000: out_v[299] = 10'b1001111111;
    16'b0000100100010000: out_v[299] = 10'b1010000100;
    16'b0000100000000000: out_v[299] = 10'b1000001010;
    16'b0000000100000001: out_v[299] = 10'b0011100111;
    16'b0000000000000000: out_v[299] = 10'b1110001100;
    16'b0000000100000000: out_v[299] = 10'b0011011101;
    16'b0000000000000001: out_v[299] = 10'b0000010101;
    16'b0000100100001001: out_v[299] = 10'b0010100011;
    16'b0000000100010001: out_v[299] = 10'b1010110111;
    16'b0000100100000001: out_v[299] = 10'b1101101100;
    16'b0000100000001000: out_v[299] = 10'b0011000011;
    16'b0000100100000000: out_v[299] = 10'b1011001100;
    16'b0000000000010001: out_v[299] = 10'b0000010111;
    16'b0000000100001001: out_v[299] = 10'b0101101010;
    16'b0000000110000001: out_v[299] = 10'b1010110011;
    16'b0000100101001001: out_v[299] = 10'b0100011001;
    16'b0000100100001000: out_v[299] = 10'b1110100001;
    16'b0010100110000001: out_v[299] = 10'b0000001100;
    16'b0000100111001101: out_v[299] = 10'b1110110011;
    16'b0010000110000001: out_v[299] = 10'b0111100100;
    16'b0010100110001000: out_v[299] = 10'b1001011000;
    16'b0000100001001101: out_v[299] = 10'b1011100100;
    16'b0000100101001000: out_v[299] = 10'b0000010100;
    16'b0010100101001001: out_v[299] = 10'b0110100110;
    16'b0000100110001001: out_v[299] = 10'b0000110101;
    16'b0010100110001001: out_v[299] = 10'b0110000100;
    16'b0010100100001001: out_v[299] = 10'b1010110111;
    16'b0000100111001000: out_v[299] = 10'b0000011110;
    16'b0000100011001001: out_v[299] = 10'b1101000110;
    16'b0000100011001101: out_v[299] = 10'b0011010011;
    16'b0010000100000000: out_v[299] = 10'b0001111011;
    16'b0000000101001000: out_v[299] = 10'b0111100100;
    16'b0010100101001000: out_v[299] = 10'b1110000111;
    16'b0000100001001100: out_v[299] = 10'b1101100101;
    16'b0010100110011001: out_v[299] = 10'b1101000101;
    16'b0000000101000001: out_v[299] = 10'b1010100100;
    16'b0010100111001001: out_v[299] = 10'b1011100001;
    16'b0010100100001000: out_v[299] = 10'b1101001011;
    16'b0000100111001001: out_v[299] = 10'b1010111011;
    16'b0000100110001000: out_v[299] = 10'b0111011001;
    16'b0000000110000000: out_v[299] = 10'b0001101011;
    16'b0000100001001001: out_v[299] = 10'b1100110011;
    16'b0010100110000000: out_v[299] = 10'b1000111111;
    16'b0010000110000000: out_v[299] = 10'b1000011100;
    16'b0000100101001101: out_v[299] = 10'b1111100111;
    16'b0000100001001000: out_v[299] = 10'b0010110010;
    16'b0010100100000000: out_v[299] = 10'b0101110110;
    16'b0010000100000001: out_v[299] = 10'b0110110100;
    16'b0000100110000000: out_v[299] = 10'b0011000111;
    16'b0000000101001001: out_v[299] = 10'b0011100101;
    16'b0000100110011001: out_v[299] = 10'b0000000101;
    16'b0000000111000001: out_v[299] = 10'b1110110101;
    16'b0000000100001000: out_v[299] = 10'b0111001100;
    16'b0010000110001000: out_v[299] = 10'b1010011101;
    16'b0000000110001000: out_v[299] = 10'b0100111010;
    16'b0010000100001000: out_v[299] = 10'b0001100011;
    16'b0001100100001001: out_v[299] = 10'b1011000011;
    16'b0010100110011000: out_v[299] = 10'b1001101001;
    16'b0000100010001000: out_v[299] = 10'b0011011010;
    16'b0000000010000000: out_v[299] = 10'b0111001100;
    16'b0010100111001000: out_v[299] = 10'b0111001000;
    16'b0001100100001000: out_v[299] = 10'b1101001001;
    16'b0000000100011000: out_v[299] = 10'b1101101000;
    16'b0011100110001000: out_v[299] = 10'b0111010111;
    16'b0010000110011000: out_v[299] = 10'b0010111001;
    16'b0000000000001000: out_v[299] = 10'b1111010000;
    16'b0000000110011000: out_v[299] = 10'b0001110100;
    16'b0010100010001000: out_v[299] = 10'b1101010101;
    16'b0000000010001000: out_v[299] = 10'b0100001011;
    16'b0000100000111001: out_v[299] = 10'b1100101111;
    16'b0000100000011001: out_v[299] = 10'b0000111100;
    16'b0010100011001000: out_v[299] = 10'b0110110001;
    16'b0000100001011001: out_v[299] = 10'b0010101011;
    16'b0010100001001001: out_v[299] = 10'b1110011010;
    16'b0010100000001000: out_v[299] = 10'b0100011011;
    16'b0000100000011000: out_v[299] = 10'b0010010011;
    16'b0000100011011000: out_v[299] = 10'b0110100011;
    16'b0000000000011001: out_v[299] = 10'b0101111001;
    16'b0010100001001000: out_v[299] = 10'b0011011110;
    16'b0010100000001001: out_v[299] = 10'b0001111101;
    16'b0000100010011000: out_v[299] = 10'b0010011111;
    16'b0000100000001001: out_v[299] = 10'b1000001111;
    16'b0010100000011001: out_v[299] = 10'b0010001011;
    16'b0000100001011000: out_v[299] = 10'b1110010010;
    16'b0000100001111001: out_v[299] = 10'b1101110110;
    16'b0000000000011000: out_v[299] = 10'b0100011101;
    16'b0000000100011001: out_v[299] = 10'b1000001001;
    16'b0000000000110011: out_v[299] = 10'b1111011111;
    16'b0000000010010000: out_v[299] = 10'b1100110011;
    16'b0000000100110010: out_v[299] = 10'b1111001110;
    16'b0000000100110011: out_v[299] = 10'b1101011110;
    16'b0000000111011000: out_v[299] = 10'b0111100010;
    16'b0000000100100011: out_v[299] = 10'b1111110101;
    16'b0010100110010000: out_v[299] = 10'b0010111110;
    16'b0000000010011000: out_v[299] = 10'b1010100010;
    16'b0000000100111011: out_v[299] = 10'b0001110101;
    16'b0000000000100011: out_v[299] = 10'b1011010101;
    16'b0010000000001000: out_v[299] = 10'b1000110111;
    16'b0010000110010000: out_v[299] = 10'b0011110000;
    16'b0000000000010000: out_v[299] = 10'b0010101100;
    16'b0000000101011000: out_v[299] = 10'b1110111010;
    16'b0000000000110010: out_v[299] = 10'b0001011011;
    16'b0000000110011100: out_v[299] = 10'b0110011111;
    16'b0000000111011101: out_v[299] = 10'b0110000011;
    16'b0000000110011101: out_v[299] = 10'b0010110011;
    16'b0010100011001001: out_v[299] = 10'b0010010100;
    16'b0000100100011101: out_v[299] = 10'b0010110111;
    16'b0010000010001001: out_v[299] = 10'b1110111001;
    16'b0000100101011101: out_v[299] = 10'b0111111011;
    16'b0000000100000100: out_v[299] = 10'b1011010011;
    16'b0000000110011001: out_v[299] = 10'b0010000011;
    16'b0000100010010001: out_v[299] = 10'b1011100100;
    16'b0000000101011101: out_v[299] = 10'b0111001010;
    16'b0000000110010100: out_v[299] = 10'b0110110101;
    16'b0010100001000001: out_v[299] = 10'b0111101001;
    16'b0000100000010001: out_v[299] = 10'b1001100010;
    16'b0010000011001001: out_v[299] = 10'b1011010010;
    16'b0000000010011001: out_v[299] = 10'b0111101111;
    16'b0000000100001101: out_v[299] = 10'b0111010001;
    16'b0000100111011101: out_v[299] = 10'b0101010111;
    16'b0000000100011101: out_v[299] = 10'b0111101011;
    16'b0000000110000100: out_v[299] = 10'b1010000101;
    16'b0010100011011001: out_v[299] = 10'b1011101111;
    16'b0000000110001100: out_v[299] = 10'b0110010001;
    16'b0000000010011100: out_v[299] = 10'b1110100110;
    16'b0000100010011001: out_v[299] = 10'b1101010011;
    16'b0000000100001100: out_v[299] = 10'b1011111001;
    16'b0010100011000001: out_v[299] = 10'b1011101010;
    16'b0000000011011001: out_v[299] = 10'b1111100101;
    16'b0000000111011100: out_v[299] = 10'b0101010111;
    16'b0000000100000101: out_v[299] = 10'b1010110110;
    16'b0000000101001101: out_v[299] = 10'b0100101111;
    16'b0000000101011001: out_v[299] = 10'b0101011110;
    16'b0000000100011100: out_v[299] = 10'b0010101110;
    16'b0000000001011001: out_v[299] = 10'b1001101110;
    16'b0000000110010101: out_v[299] = 10'b0101011111;
    16'b0000100010010000: out_v[299] = 10'b1000110010;
    16'b0000000010011101: out_v[299] = 10'b0100111111;
    16'b0000100011011001: out_v[299] = 10'b0010111101;
    16'b0010100010000001: out_v[299] = 10'b0011100000;
    16'b0010100000011000: out_v[299] = 10'b0110100011;
    16'b0010100100011001: out_v[299] = 10'b1011000111;
    16'b0010100100011000: out_v[299] = 10'b1101110011;
    16'b0010100010011000: out_v[299] = 10'b1000111010;
    16'b0010100000010000: out_v[299] = 10'b0111100001;
    16'b0010100010010000: out_v[299] = 10'b0110110011;
    16'b0010100100000001: out_v[299] = 10'b1100111011;
    16'b0000100000010000: out_v[299] = 10'b0101110000;
    16'b0010000100001001: out_v[299] = 10'b1000000111;
    16'b0000100100010001: out_v[299] = 10'b1101001001;
    16'b0000100100111011: out_v[299] = 10'b0101011101;
    16'b0000100100111010: out_v[299] = 10'b0011010011;
    16'b0000100100111001: out_v[299] = 10'b0001101110;
    16'b0010100111011000: out_v[299] = 10'b1100000010;
    16'b0000100100111000: out_v[299] = 10'b0010010110;
    16'b0000100100110001: out_v[299] = 10'b0111010110;
    default: out_v[299] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000101000000: out_v[300] = 10'b1000110000;
    16'b0110000111000001: out_v[300] = 10'b0000101111;
    16'b0110000111000000: out_v[300] = 10'b0010110110;
    16'b0110000101000000: out_v[300] = 10'b0010101101;
    16'b0110000101000001: out_v[300] = 10'b1100100011;
    16'b0100000001000000: out_v[300] = 10'b0010001010;
    16'b0010000110000000: out_v[300] = 10'b1011000011;
    16'b0110000100000000: out_v[300] = 10'b0101000100;
    16'b0110000110000000: out_v[300] = 10'b0001001100;
    16'b0010000111000000: out_v[300] = 10'b0010110100;
    16'b0010000101000000: out_v[300] = 10'b0010001111;
    16'b0110000110000001: out_v[300] = 10'b0101000010;
    16'b0100000001000001: out_v[300] = 10'b1111000001;
    16'b0111000110000000: out_v[300] = 10'b1000001011;
    16'b0000000011000000: out_v[300] = 10'b0011100011;
    16'b0010000101000001: out_v[300] = 10'b1100010011;
    16'b0110000011000001: out_v[300] = 10'b0001111011;
    16'b0110000001000000: out_v[300] = 10'b0110010000;
    16'b0000000001000000: out_v[300] = 10'b1000011001;
    16'b0010000111000001: out_v[300] = 10'b0010101001;
    16'b0110000101110000: out_v[300] = 10'b0000101001;
    16'b0111000111000000: out_v[300] = 10'b1010111111;
    16'b0111000111000001: out_v[300] = 10'b1101011011;
    16'b0100000011000001: out_v[300] = 10'b0001011010;
    16'b0010000100000000: out_v[300] = 10'b1110110111;
    16'b0010000100000001: out_v[300] = 10'b0110111110;
    16'b0110000000000001: out_v[300] = 10'b0110110100;
    16'b0110000100000001: out_v[300] = 10'b0001111010;
    16'b0000000011000001: out_v[300] = 10'b1000111111;
    16'b0100000000000001: out_v[300] = 10'b0110110010;
    16'b0110000001000001: out_v[300] = 10'b1101001011;
    16'b0110000000000000: out_v[300] = 10'b1001110100;
    16'b0100000011000000: out_v[300] = 10'b0010110010;
    16'b0100000000000000: out_v[300] = 10'b0111010001;
    16'b0000000100000001: out_v[300] = 10'b1000011010;
    16'b0010000000000000: out_v[300] = 10'b1100010111;
    16'b0010000000000001: out_v[300] = 10'b1100000101;
    16'b0100101001000000: out_v[300] = 10'b0110001111;
    16'b0110000100110000: out_v[300] = 10'b0001100101;
    16'b0100100001000000: out_v[300] = 10'b0100110110;
    16'b0100000001110000: out_v[300] = 10'b0101000110;
    16'b0110000011000000: out_v[300] = 10'b0010101001;
    16'b0010000101110000: out_v[300] = 10'b1100100010;
    16'b0110101110000000: out_v[300] = 10'b1100100111;
    16'b0100000010000000: out_v[300] = 10'b1011101111;
    16'b0100101011000000: out_v[300] = 10'b0111111111;
    16'b0110000101110001: out_v[300] = 10'b1111000000;
    16'b0110000010000000: out_v[300] = 10'b1101001110;
    16'b0100101010000000: out_v[300] = 10'b0110011101;
    16'b0000000001000001: out_v[300] = 10'b0111001011;
    16'b0110000100110001: out_v[300] = 10'b1010101010;
    16'b0110101101000000: out_v[300] = 10'b0100000011;
    16'b0110101111000000: out_v[300] = 10'b0101100101;
    16'b0110100101000000: out_v[300] = 10'b0110000111;
    16'b0000000000000001: out_v[300] = 10'b1010101111;
    16'b0100000000110000: out_v[300] = 10'b1101100111;
    16'b0000000000000000: out_v[300] = 10'b1001111111;
    16'b0110000111110000: out_v[300] = 10'b0010010011;
    16'b0000000010000000: out_v[300] = 10'b0110010010;
    16'b0110000001110000: out_v[300] = 10'b1111110011;
    16'b0110100101000001: out_v[300] = 10'b0000001111;
    16'b0000000101000001: out_v[300] = 10'b0110011001;
    16'b0110101111000001: out_v[300] = 10'b0010001010;
    16'b0000000000110001: out_v[300] = 10'b0011011010;
    16'b0010000101110001: out_v[300] = 10'b0011001010;
    16'b0000000101110001: out_v[300] = 10'b0111010001;
    16'b0000000001110000: out_v[300] = 10'b0010011010;
    16'b0000000100110001: out_v[300] = 10'b1000110111;
    16'b0010000100110001: out_v[300] = 10'b0111011101;
    16'b0000000001110001: out_v[300] = 10'b0000111010;
    16'b0110000111110001: out_v[300] = 10'b0101001101;
    16'b0010000111110001: out_v[300] = 10'b0100110010;
    16'b0010000110000001: out_v[300] = 10'b1010110010;
    16'b0000000000110000: out_v[300] = 10'b0010011001;
    16'b0000000100000000: out_v[300] = 10'b0010110001;
    16'b0000000111000000: out_v[300] = 10'b0101010111;
    16'b0000000110000000: out_v[300] = 10'b1100101010;
    16'b0000000011110000: out_v[300] = 10'b0110100011;
    16'b0101000000000001: out_v[300] = 10'b1010100011;
    16'b0111000101000001: out_v[300] = 10'b1011110110;
    16'b0000000111000001: out_v[300] = 10'b0101110101;
    16'b0110101100000001: out_v[300] = 10'b1101000000;
    16'b0000000010000001: out_v[300] = 10'b1001100111;
    16'b0000000110000001: out_v[300] = 10'b1101000011;
    16'b0110101100000000: out_v[300] = 10'b0001111010;
    16'b0110100100000001: out_v[300] = 10'b1001101100;
    16'b0110001100000000: out_v[300] = 10'b0011111001;
    16'b0110100100000000: out_v[300] = 10'b1011010011;
    16'b0110001100000001: out_v[300] = 10'b1010000111;
    16'b0100101000000001: out_v[300] = 10'b1111101011;
    16'b0110101000000001: out_v[300] = 10'b1111100000;
    16'b0110101000000000: out_v[300] = 10'b1000111011;
    16'b0100101000000000: out_v[300] = 10'b0011000001;
    16'b0110001101000001: out_v[300] = 10'b0110110001;
    16'b0110101101000001: out_v[300] = 10'b0101011011;
    16'b0010000100110000: out_v[300] = 10'b0110000010;
    16'b0010000001000000: out_v[300] = 10'b0110011001;
    16'b0000000101110000: out_v[300] = 10'b1111000111;
    16'b0110000010000001: out_v[300] = 10'b1010000111;
    16'b0100000101000000: out_v[300] = 10'b1101111010;
    16'b0100000101000001: out_v[300] = 10'b1111010010;
    default: out_v[300] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000100010100000: out_v[301] = 10'b0101011000;
    16'b1000100010000000: out_v[301] = 10'b1111001001;
    16'b1000000011000000: out_v[301] = 10'b0011000111;
    16'b1000000011100000: out_v[301] = 10'b0010111111;
    16'b1000100000100000: out_v[301] = 10'b0111011001;
    16'b1000100010101000: out_v[301] = 10'b1001010001;
    16'b1000000010000000: out_v[301] = 10'b0010110110;
    16'b1000000000000000: out_v[301] = 10'b1110011001;
    16'b0000000010000000: out_v[301] = 10'b0101100011;
    16'b1000000001000000: out_v[301] = 10'b1111001011;
    16'b1000100011100000: out_v[301] = 10'b1010001001;
    16'b0000100000100000: out_v[301] = 10'b1110111001;
    16'b1100000001000000: out_v[301] = 10'b0011001001;
    16'b1000100001100000: out_v[301] = 10'b1011011000;
    16'b1000100000000000: out_v[301] = 10'b0100101101;
    16'b1000000010001000: out_v[301] = 10'b0011110011;
    16'b0000100010101000: out_v[301] = 10'b0000111011;
    16'b1100100011100000: out_v[301] = 10'b0101100100;
    16'b1000100000101000: out_v[301] = 10'b1000011001;
    16'b0000000001000000: out_v[301] = 10'b0000010101;
    16'b1100000011000000: out_v[301] = 10'b1011001001;
    16'b1000100010100000: out_v[301] = 10'b1111010110;
    16'b1100100001100000: out_v[301] = 10'b0011110000;
    16'b0100000001000000: out_v[301] = 10'b1010111011;
    16'b0000000011000000: out_v[301] = 10'b0010110110;
    16'b1000100010001000: out_v[301] = 10'b0000011111;
    16'b0000100000101000: out_v[301] = 10'b1110010110;
    16'b1000100011101000: out_v[301] = 10'b0001011011;
    16'b0000000000000000: out_v[301] = 10'b1010111011;
    16'b0000000010001000: out_v[301] = 10'b0110111100;
    16'b0100000010000000: out_v[301] = 10'b0000010110;
    16'b0100000011000000: out_v[301] = 10'b0110000101;
    16'b0100000000000000: out_v[301] = 10'b1000100110;
    16'b0000000000001000: out_v[301] = 10'b0100110001;
    16'b0100100000101000: out_v[301] = 10'b0101010110;
    16'b0000100001101000: out_v[301] = 10'b1110100101;
    16'b0100000000001000: out_v[301] = 10'b1110100011;
    16'b0000000001001000: out_v[301] = 10'b1001010110;
    16'b0000100011101000: out_v[301] = 10'b0011011110;
    16'b0100100000100000: out_v[301] = 10'b0000110111;
    16'b0000000011001000: out_v[301] = 10'b0010010110;
    16'b0100100001101000: out_v[301] = 10'b1000011011;
    16'b0000000001101000: out_v[301] = 10'b1101100110;
    16'b1000100001101000: out_v[301] = 10'b0001000110;
    16'b0000000000101000: out_v[301] = 10'b1101011101;
    16'b0000100001100000: out_v[301] = 10'b0111101011;
    16'b0100000001001000: out_v[301] = 10'b0110111011;
    16'b0000000000100000: out_v[301] = 10'b0101011110;
    16'b0000000001100000: out_v[301] = 10'b1101100010;
    16'b0000100000000000: out_v[301] = 10'b0110110101;
    16'b0100100010101000: out_v[301] = 10'b1000010100;
    16'b0100000000100000: out_v[301] = 10'b1001110111;
    16'b0000100011000000: out_v[301] = 10'b0001011010;
    16'b0000000000001001: out_v[301] = 10'b0001111111;
    16'b0000100000001000: out_v[301] = 10'b1101100010;
    16'b0000100010000000: out_v[301] = 10'b0110100001;
    16'b0100100001100000: out_v[301] = 10'b1011111000;
    16'b0100000010001000: out_v[301] = 10'b0111000001;
    16'b0100101011100000: out_v[301] = 10'b1100001111;
    16'b0000000010101000: out_v[301] = 10'b0101001010;
    16'b0000000000000001: out_v[301] = 10'b1001011011;
    16'b0000100010001000: out_v[301] = 10'b0010101011;
    16'b0000100011100000: out_v[301] = 10'b1100110010;
    16'b0100100011100000: out_v[301] = 10'b0111011011;
    16'b1000000000001000: out_v[301] = 10'b0100101111;
    16'b0100000011001000: out_v[301] = 10'b0101001010;
    16'b0100100001000000: out_v[301] = 10'b1111000010;
    16'b1100100011000000: out_v[301] = 10'b0110110110;
    16'b0100100011000000: out_v[301] = 10'b1101011001;
    16'b0000100001000000: out_v[301] = 10'b1100110001;
    16'b0000000010001001: out_v[301] = 10'b0101110001;
    16'b0000000010000001: out_v[301] = 10'b1101001001;
    16'b1000100000001000: out_v[301] = 10'b1101001110;
    16'b1100100000101000: out_v[301] = 10'b0000011110;
    16'b1000100000101001: out_v[301] = 10'b0011011111;
    16'b1000000000100000: out_v[301] = 10'b0100010101;
    16'b1000100010101001: out_v[301] = 10'b1111000000;
    16'b1000100000100001: out_v[301] = 10'b0010111110;
    16'b1000000000101000: out_v[301] = 10'b1011001110;
    16'b1000000010100000: out_v[301] = 10'b1100101000;
    16'b1100100000100000: out_v[301] = 10'b1100101010;
    16'b1100100001101000: out_v[301] = 10'b0110010100;
    16'b1000000010000001: out_v[301] = 10'b1100100111;
    16'b1000000010001001: out_v[301] = 10'b1000111110;
    16'b1100100001000000: out_v[301] = 10'b0011001001;
    16'b1000100001000000: out_v[301] = 10'b1111111010;
    16'b1000000001100000: out_v[301] = 10'b1100101110;
    16'b0001100010100001: out_v[301] = 10'b0101111111;
    16'b0000101010101000: out_v[301] = 10'b0100100110;
    16'b0001000010000001: out_v[301] = 10'b0111101101;
    16'b0000000010100000: out_v[301] = 10'b0110011001;
    16'b1001000010000001: out_v[301] = 10'b1001100000;
    16'b1001100010101001: out_v[301] = 10'b1000000001;
    16'b0000100010101001: out_v[301] = 10'b1111100010;
    16'b0000001010001000: out_v[301] = 10'b1011110011;
    16'b1001000010100001: out_v[301] = 10'b1001001110;
    16'b1001100010100001: out_v[301] = 10'b0111000111;
    16'b0000101010101001: out_v[301] = 10'b0111110001;
    16'b0001000010100001: out_v[301] = 10'b1100111111;
    16'b0000100010100001: out_v[301] = 10'b0111100100;
    16'b0001101010101001: out_v[301] = 10'b1100111000;
    16'b0001100010101001: out_v[301] = 10'b1101010111;
    16'b0000101010100000: out_v[301] = 10'b1110100101;
    16'b0000000010100001: out_v[301] = 10'b0001111111;
    16'b0000001010000000: out_v[301] = 10'b0101011010;
    16'b1000101010101000: out_v[301] = 10'b0111100011;
    16'b1000100010100001: out_v[301] = 10'b1101101111;
    16'b1000000010101000: out_v[301] = 10'b0111100000;
    16'b1100000010001000: out_v[301] = 10'b1101010111;
    16'b1000000000100001: out_v[301] = 10'b1001110110;
    16'b1000000010100001: out_v[301] = 10'b1111101000;
    16'b1100100010101000: out_v[301] = 10'b0010110111;
    16'b1000000000000001: out_v[301] = 10'b1010101110;
    default: out_v[301] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000010111010001: out_v[302] = 10'b1001101010;
    16'b0000011110010001: out_v[302] = 10'b1001100101;
    16'b0001011111010001: out_v[302] = 10'b0101100011;
    16'b0001011110010001: out_v[302] = 10'b0100000000;
    16'b0000010101010001: out_v[302] = 10'b0110001011;
    16'b0000010010010001: out_v[302] = 10'b1100101011;
    16'b0001010010010001: out_v[302] = 10'b0100011001;
    16'b0000011101000001: out_v[302] = 10'b1111000111;
    16'b0001001110010001: out_v[302] = 10'b1011000010;
    16'b0000010110010001: out_v[302] = 10'b0000110011;
    16'b0000011111010001: out_v[302] = 10'b1011100000;
    16'b0000011111000001: out_v[302] = 10'b0110000001;
    16'b0000011101010001: out_v[302] = 10'b0001011110;
    16'b0001011010010001: out_v[302] = 10'b0000111111;
    16'b0001011100010001: out_v[302] = 10'b0110111010;
    16'b0001010010000001: out_v[302] = 10'b1111111011;
    16'b0001011110000001: out_v[302] = 10'b1101100110;
    16'b0000011011000001: out_v[302] = 10'b0101110011;
    16'b0000010010000001: out_v[302] = 10'b1110100001;
    16'b0000010000010001: out_v[302] = 10'b1001010011;
    16'b0001001110010000: out_v[302] = 10'b0111111001;
    16'b0001010110010001: out_v[302] = 10'b1010001101;
    16'b0000010100010001: out_v[302] = 10'b0111011011;
    16'b0001011111000001: out_v[302] = 10'b0011001111;
    16'b0000000010000001: out_v[302] = 10'b1110001000;
    16'b0000011001000001: out_v[302] = 10'b1111001111;
    16'b0000010000000001: out_v[302] = 10'b1001001011;
    16'b0000011100010001: out_v[302] = 10'b1011111011;
    16'b0001011101000001: out_v[302] = 10'b0110000101;
    16'b0000011110000001: out_v[302] = 10'b1010111100;
    16'b0001011100000001: out_v[302] = 10'b1110001010;
    16'b0000011100000001: out_v[302] = 10'b1100000111;
    16'b0000000010000000: out_v[302] = 10'b1011001100;
    16'b0000000011000000: out_v[302] = 10'b1001110010;
    16'b0000000000000001: out_v[302] = 10'b0001110011;
    16'b0000000001000000: out_v[302] = 10'b1100110101;
    16'b0000000000000000: out_v[302] = 10'b1010100000;
    16'b0000010000000000: out_v[302] = 10'b0110011101;
    16'b0000000110000000: out_v[302] = 10'b1000010010;
    16'b0000000011100000: out_v[302] = 10'b0100011101;
    16'b0000011000010001: out_v[302] = 10'b0110111011;
    16'b0000010100000001: out_v[302] = 10'b0011010100;
    16'b0000010110000001: out_v[302] = 10'b1001110110;
    16'b0000000100000001: out_v[302] = 10'b1011001111;
    16'b0001011000010001: out_v[302] = 10'b1111101110;
    16'b0000010001000001: out_v[302] = 10'b0000010110;
    16'b0000001010010000: out_v[302] = 10'b0000011101;
    16'b0001010100010001: out_v[302] = 10'b1101011110;
    16'b0000010100100001: out_v[302] = 10'b0010001011;
    16'b0001010100000001: out_v[302] = 10'b1111110101;
    16'b0001010110000001: out_v[302] = 10'b0101000110;
    16'b0001010100000000: out_v[302] = 10'b0011101110;
    16'b0001010000000001: out_v[302] = 10'b1111111000;
    16'b0000010011000001: out_v[302] = 10'b0100101100;
    16'b0000000110100000: out_v[302] = 10'b1100010100;
    16'b0000010000100001: out_v[302] = 10'b1111101011;
    16'b0000000100000000: out_v[302] = 10'b0010101110;
    16'b0000010001100001: out_v[302] = 10'b1000001100;
    16'b0000000010100000: out_v[302] = 10'b0111010001;
    16'b0000010011100001: out_v[302] = 10'b0010100111;
    16'b0010001010010000: out_v[302] = 10'b1100101101;
    16'b0000001110010000: out_v[302] = 10'b0101100101;
    16'b0000000101010001: out_v[302] = 10'b0001001010;
    16'b0000001011110000: out_v[302] = 10'b0111001001;
    16'b0000000111100000: out_v[302] = 10'b0011101001;
    16'b0000001111110001: out_v[302] = 10'b1011000111;
    16'b0000010111000001: out_v[302] = 10'b1101000001;
    16'b0000000111000000: out_v[302] = 10'b1010011001;
    16'b0000000111010001: out_v[302] = 10'b0000110001;
    16'b0000000111110000: out_v[302] = 10'b1001001111;
    16'b0000000111010000: out_v[302] = 10'b1101101001;
    16'b0000001011100000: out_v[302] = 10'b0111011011;
    16'b0000001111100000: out_v[302] = 10'b1101011111;
    16'b0000000101010000: out_v[302] = 10'b0001100100;
    16'b0000011111110001: out_v[302] = 10'b0100100111;
    16'b0000010101110001: out_v[302] = 10'b1111011111;
    16'b0000010101100001: out_v[302] = 10'b0011011011;
    16'b0000011101110001: out_v[302] = 10'b0110111011;
    16'b0000000110010000: out_v[302] = 10'b0101011010;
    16'b0000011101100001: out_v[302] = 10'b1010111011;
    16'b0001010101010001: out_v[302] = 10'b1111110111;
    16'b0000000100010001: out_v[302] = 10'b1101011101;
    16'b0000001111110000: out_v[302] = 10'b1011011010;
    16'b0000000001000001: out_v[302] = 10'b1101010110;
    16'b0000001101110001: out_v[302] = 10'b0111110011;
    16'b0000001111010000: out_v[302] = 10'b1101001110;
    16'b0000000011000001: out_v[302] = 10'b1111100100;
    16'b0000010101000001: out_v[302] = 10'b1111011001;
    16'b0000010111110001: out_v[302] = 10'b1011110111;
    16'b0000000101110001: out_v[302] = 10'b1110100010;
    16'b0000010010000000: out_v[302] = 10'b0110110000;
    16'b0000010001000000: out_v[302] = 10'b0011100111;
    16'b0000010100110001: out_v[302] = 10'b0100011001;
    16'b0001010000000000: out_v[302] = 10'b1110101001;
    16'b0000000100010000: out_v[302] = 10'b0101110001;
    16'b0000001111010001: out_v[302] = 10'b0010111111;
    16'b0000001111000001: out_v[302] = 10'b0110110011;
    16'b0000000111000001: out_v[302] = 10'b0111111111;
    16'b0000001101010000: out_v[302] = 10'b0010110111;
    16'b0001010010000000: out_v[302] = 10'b0001110011;
    16'b0000001001000000: out_v[302] = 10'b0110100000;
    16'b0000001100010000: out_v[302] = 10'b0010110010;
    16'b0000001101000000: out_v[302] = 10'b1111110110;
    16'b0000000110010001: out_v[302] = 10'b1110100101;
    16'b0000001101010001: out_v[302] = 10'b1011011110;
    16'b0001000000000000: out_v[302] = 10'b0001100110;
    16'b0000000010010000: out_v[302] = 10'b1001001001;
    16'b0000001100000000: out_v[302] = 10'b0011000010;
    16'b0000000010010001: out_v[302] = 10'b0101100010;
    16'b0000000000010000: out_v[302] = 10'b0011001001;
    16'b0000001100110000: out_v[302] = 10'b0101100000;
    16'b0000001000010000: out_v[302] = 10'b1011000111;
    16'b0000001110000000: out_v[302] = 10'b1011011111;
    16'b0000001000000000: out_v[302] = 10'b1011011011;
    16'b0000001110010001: out_v[302] = 10'b0110001111;
    16'b0000001100100000: out_v[302] = 10'b0101101011;
    16'b0000010010100001: out_v[302] = 10'b1010010111;
    16'b0000010010000100: out_v[302] = 10'b0001111011;
    16'b0000010011000101: out_v[302] = 10'b1000111101;
    16'b0000010011000000: out_v[302] = 10'b0001111110;
    16'b0000000011000100: out_v[302] = 10'b0111110011;
    16'b0000010010000101: out_v[302] = 10'b0110001101;
    16'b0000010011000100: out_v[302] = 10'b0010100111;
    16'b0000010111010100: out_v[302] = 10'b0111111111;
    16'b0000000101000000: out_v[302] = 10'b0110101011;
    16'b0000000101000001: out_v[302] = 10'b1111011011;
    16'b0000010011010001: out_v[302] = 10'b0011100111;
    default: out_v[302] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001000001100100: out_v[303] = 10'b0011111011;
    16'b1000000100100100: out_v[303] = 10'b1100000111;
    16'b0000000101100101: out_v[303] = 10'b0001010001;
    16'b0000000001100100: out_v[303] = 10'b1001001000;
    16'b1000000000100100: out_v[303] = 10'b1100001110;
    16'b1000000101100100: out_v[303] = 10'b0001001010;
    16'b0000000101100000: out_v[303] = 10'b0000001011;
    16'b0000000100100100: out_v[303] = 10'b0111011011;
    16'b0000000100100000: out_v[303] = 10'b0010111011;
    16'b1000000001100100: out_v[303] = 10'b0010010111;
    16'b0000000001100101: out_v[303] = 10'b0110100001;
    16'b1000000100100000: out_v[303] = 10'b1000011011;
    16'b1000000001100000: out_v[303] = 10'b1001110110;
    16'b1000000101100101: out_v[303] = 10'b0110000001;
    16'b0000000101000101: out_v[303] = 10'b1100001010;
    16'b0000000101100001: out_v[303] = 10'b1110100101;
    16'b0000000101100100: out_v[303] = 10'b0011011010;
    16'b0000000000100000: out_v[303] = 10'b0010011011;
    16'b0000000000100100: out_v[303] = 10'b0011011100;
    16'b1000000000000100: out_v[303] = 10'b0101000101;
    16'b0001000001100101: out_v[303] = 10'b0101100000;
    16'b0000000101000001: out_v[303] = 10'b1000111101;
    16'b1000000000100000: out_v[303] = 10'b1111011000;
    16'b0000000100000101: out_v[303] = 10'b1001011011;
    16'b1000000101000101: out_v[303] = 10'b0000110111;
    16'b0000000000000100: out_v[303] = 10'b1000100111;
    16'b1000000001100101: out_v[303] = 10'b0111100111;
    16'b0000000001100000: out_v[303] = 10'b1110011000;
    16'b0001000101100101: out_v[303] = 10'b0101100111;
    16'b0000000001000101: out_v[303] = 10'b0011001101;
    16'b1000000001000100: out_v[303] = 10'b0100010100;
    16'b1000000101100000: out_v[303] = 10'b1001111001;
    16'b0000000001000100: out_v[303] = 10'b1010100110;
    16'b0000000001100001: out_v[303] = 10'b0100100011;
    16'b0000000000000000: out_v[303] = 10'b0100011011;
    16'b1000000000000000: out_v[303] = 10'b1001100110;
    16'b0000000001000000: out_v[303] = 10'b0010001001;
    16'b1000000001000000: out_v[303] = 10'b0010101110;
    16'b1001000001000000: out_v[303] = 10'b0011100000;
    16'b1001000000000000: out_v[303] = 10'b1111100001;
    16'b1000000001000001: out_v[303] = 10'b1110000101;
    16'b1000000101000100: out_v[303] = 10'b0110011110;
    16'b1000000000000101: out_v[303] = 10'b0010110110;
    16'b1000000001000101: out_v[303] = 10'b1010000110;
    16'b0001000001000001: out_v[303] = 10'b0001011011;
    16'b0001000001000100: out_v[303] = 10'b0111000110;
    16'b0001000001000000: out_v[303] = 10'b0000011101;
    16'b0001000001100000: out_v[303] = 10'b1011101110;
    16'b0000000001000001: out_v[303] = 10'b1001001000;
    16'b0001000001100001: out_v[303] = 10'b1010100110;
    16'b1000000000100001: out_v[303] = 10'b0011010010;
    16'b1000000000000001: out_v[303] = 10'b0101110011;
    16'b1001000001100001: out_v[303] = 10'b1101101011;
    16'b1001000000100000: out_v[303] = 10'b0101011111;
    16'b0000000000100001: out_v[303] = 10'b1110010010;
    16'b1001000001100000: out_v[303] = 10'b1100000110;
    16'b1000000001100001: out_v[303] = 10'b1101100110;
    16'b0000000000000001: out_v[303] = 10'b0010111001;
    16'b1001000000100001: out_v[303] = 10'b0101111111;
    16'b1000000000100101: out_v[303] = 10'b0110110010;
    16'b1000000010100000: out_v[303] = 10'b0111101110;
    16'b0000000000100101: out_v[303] = 10'b1110010100;
    16'b1000000010100100: out_v[303] = 10'b1000101110;
    16'b1000000100100101: out_v[303] = 10'b0111110010;
    16'b1000000100000101: out_v[303] = 10'b0001010011;
    16'b0001000000100001: out_v[303] = 10'b0111000011;
    16'b1001000000000001: out_v[303] = 10'b0010110000;
    16'b1001000001000001: out_v[303] = 10'b1000011011;
    16'b0001000000000001: out_v[303] = 10'b1111101101;
    16'b1001000001100101: out_v[303] = 10'b0011011010;
    16'b1001000001100100: out_v[303] = 10'b1110100010;
    16'b1001000001000100: out_v[303] = 10'b0101111100;
    16'b0000100001100001: out_v[303] = 10'b1001100010;
    16'b1000100001000001: out_v[303] = 10'b1011001001;
    16'b0000100001000001: out_v[303] = 10'b1111001111;
    default: out_v[303] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000000010000: out_v[304] = 10'b0100101011;
    16'b0100000001010000: out_v[304] = 10'b0001000011;
    16'b0100010000010000: out_v[304] = 10'b0001110000;
    16'b0100010000000000: out_v[304] = 10'b0101001100;
    16'b0100000000010000: out_v[304] = 10'b0100001101;
    16'b0100000000000000: out_v[304] = 10'b0111011000;
    16'b0000000001010001: out_v[304] = 10'b0100101010;
    16'b0000010000000000: out_v[304] = 10'b1001001111;
    16'b0100010001010001: out_v[304] = 10'b0100110011;
    16'b0000010000010000: out_v[304] = 10'b0100010100;
    16'b0100000001010001: out_v[304] = 10'b0100000001;
    16'b0100010001010000: out_v[304] = 10'b0111010011;
    16'b0100010001000000: out_v[304] = 10'b0001011011;
    16'b0000000000000000: out_v[304] = 10'b1000111010;
    16'b0100010001000001: out_v[304] = 10'b1001110001;
    16'b0100000001000001: out_v[304] = 10'b0011110000;
    16'b0000010001000000: out_v[304] = 10'b0010001101;
    16'b0000010001000001: out_v[304] = 10'b0111000010;
    16'b0001010000010000: out_v[304] = 10'b0100001100;
    16'b0000010001010001: out_v[304] = 10'b0100000100;
    16'b0001010000000000: out_v[304] = 10'b0010001111;
    16'b0000010001010000: out_v[304] = 10'b0000101010;
    16'b0000010000010001: out_v[304] = 10'b1001101100;
    16'b0001010001000001: out_v[304] = 10'b0011110101;
    16'b0001010001010001: out_v[304] = 10'b1101001010;
    16'b0000010000000001: out_v[304] = 10'b0011100101;
    16'b1000010000000000: out_v[304] = 10'b1110001111;
    16'b0000000000010001: out_v[304] = 10'b0100001110;
    16'b0010000000000000: out_v[304] = 10'b0010010011;
    16'b0000000001000001: out_v[304] = 10'b0110011100;
    16'b0000000001010000: out_v[304] = 10'b0000011110;
    16'b0010000001000001: out_v[304] = 10'b0011011110;
    16'b0000000000000001: out_v[304] = 10'b0111110001;
    16'b0000000001000000: out_v[304] = 10'b1110011100;
    16'b0010000001010001: out_v[304] = 10'b1101010010;
    16'b0110010000010000: out_v[304] = 10'b1011101110;
    16'b0100000000000001: out_v[304] = 10'b0001111111;
    16'b0010010000010000: out_v[304] = 10'b0111010001;
    16'b0100000001000000: out_v[304] = 10'b0111110010;
    16'b0010010000000000: out_v[304] = 10'b0000111010;
    16'b0010000000010000: out_v[304] = 10'b0101100111;
    16'b1000000000000000: out_v[304] = 10'b1011011100;
    16'b1100010000000000: out_v[304] = 10'b1110110110;
    16'b0010010001110000: out_v[304] = 10'b0010111111;
    16'b0010010001010000: out_v[304] = 10'b1111000011;
    16'b0010010000110000: out_v[304] = 10'b0110000101;
    16'b0010010001010001: out_v[304] = 10'b1011001010;
    16'b0010010000010001: out_v[304] = 10'b1100100101;
    16'b0010000001000000: out_v[304] = 10'b0011101000;
    16'b0010000000110000: out_v[304] = 10'b1001000110;
    16'b0010000001110001: out_v[304] = 10'b0101111101;
    16'b0010010001110001: out_v[304] = 10'b0001111011;
    16'b0110000000000000: out_v[304] = 10'b1111000011;
    16'b0010000001010000: out_v[304] = 10'b0000111111;
    16'b0010010001000001: out_v[304] = 10'b0001101101;
    16'b0010000001110000: out_v[304] = 10'b0111110011;
    16'b0110000000010000: out_v[304] = 10'b1010100010;
    default: out_v[304] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000101000000001: out_v[305] = 10'b1010100101;
    16'b0001101000010001: out_v[305] = 10'b1100010110;
    16'b0000100000000000: out_v[305] = 10'b0110011100;
    16'b0000101000000000: out_v[305] = 10'b0011001101;
    16'b0001101000000000: out_v[305] = 10'b0001011001;
    16'b0001101000000001: out_v[305] = 10'b1010111100;
    16'b0001101010000000: out_v[305] = 10'b0011001011;
    16'b0001101000000100: out_v[305] = 10'b1111011110;
    16'b0000101010000001: out_v[305] = 10'b0001001110;
    16'b0001000000000001: out_v[305] = 10'b1101001011;
    16'b0000100000000001: out_v[305] = 10'b0101110110;
    16'b0000000000000000: out_v[305] = 10'b1101110011;
    16'b0001101000010000: out_v[305] = 10'b1101011001;
    16'b0011000000010000: out_v[305] = 10'b1100010011;
    16'b0111000000010001: out_v[305] = 10'b0100010111;
    16'b0000000000010000: out_v[305] = 10'b1100001010;
    16'b0001101000000101: out_v[305] = 10'b1110100110;
    16'b0011101000010000: out_v[305] = 10'b0011111111;
    16'b0000101010000000: out_v[305] = 10'b1001101110;
    16'b0011001000010000: out_v[305] = 10'b0101011011;
    16'b0001101010000001: out_v[305] = 10'b0010110111;
    16'b0001101010000101: out_v[305] = 10'b0001110011;
    16'b0000001000000001: out_v[305] = 10'b0101111001;
    16'b0000001000000000: out_v[305] = 10'b1101011100;
    16'b0100000000000000: out_v[305] = 10'b0001101101;
    16'b0000101000000101: out_v[305] = 10'b0101000000;
    16'b0000101000010000: out_v[305] = 10'b0111001110;
    16'b0000000000000001: out_v[305] = 10'b0111001001;
    16'b0111000000010000: out_v[305] = 10'b1010100001;
    16'b0001000000000000: out_v[305] = 10'b0111100110;
    16'b0001001000010000: out_v[305] = 10'b0111011001;
    16'b0001101010010000: out_v[305] = 10'b1111000000;
    16'b0000000010000001: out_v[305] = 10'b0010100011;
    16'b0000001010000000: out_v[305] = 10'b0100000000;
    16'b0000000010000000: out_v[305] = 10'b1010110101;
    16'b0100001010000000: out_v[305] = 10'b1011010011;
    16'b0100001000000000: out_v[305] = 10'b0100010110;
    16'b0000001010000001: out_v[305] = 10'b0011100010;
    16'b0010101010000000: out_v[305] = 10'b0100010111;
    16'b0010101000000000: out_v[305] = 10'b1101011111;
    16'b0010001010000001: out_v[305] = 10'b0111010101;
    16'b0010101010000001: out_v[305] = 10'b1000010001;
    16'b0000100010000000: out_v[305] = 10'b1110000100;
    16'b0010101010010000: out_v[305] = 10'b0101110111;
    16'b0000101010010000: out_v[305] = 10'b1101011011;
    16'b0010000010000000: out_v[305] = 10'b0011000100;
    16'b0010000000000000: out_v[305] = 10'b1001011000;
    16'b0000101000010001: out_v[305] = 10'b1011110111;
    16'b0000110000000100: out_v[305] = 10'b1010100111;
    16'b0000101000000100: out_v[305] = 10'b0000111111;
    16'b0010100010000000: out_v[305] = 10'b1110001101;
    16'b0010100000000100: out_v[305] = 10'b1011111000;
    16'b0010101010010001: out_v[305] = 10'b0110101100;
    16'b0010100000000000: out_v[305] = 10'b0011000101;
    16'b0010101000010001: out_v[305] = 10'b0001010110;
    16'b0000010000000100: out_v[305] = 10'b1000011101;
    16'b0010101000010000: out_v[305] = 10'b0011101110;
    16'b0010001010000000: out_v[305] = 10'b1010011111;
    16'b0010001000000000: out_v[305] = 10'b0110001001;
    16'b0000000000000100: out_v[305] = 10'b0001110111;
    16'b0010001010010000: out_v[305] = 10'b0101101011;
    16'b0000111000000100: out_v[305] = 10'b1100000101;
    16'b0010000000000100: out_v[305] = 10'b1010010110;
    16'b0010101000000100: out_v[305] = 10'b0100000111;
    16'b0010000010010000: out_v[305] = 10'b1100111010;
    16'b0010101000000001: out_v[305] = 10'b0110100110;
    16'b0000100000000100: out_v[305] = 10'b0011100110;
    16'b0000001000000100: out_v[305] = 10'b0011100110;
    16'b0100100010010001: out_v[305] = 10'b0111110111;
    16'b0100000000000001: out_v[305] = 10'b1101010111;
    16'b0000111010000101: out_v[305] = 10'b1001110100;
    16'b0000101010000100: out_v[305] = 10'b1000111010;
    16'b0100100010000001: out_v[305] = 10'b1101111000;
    16'b0100000010000000: out_v[305] = 10'b0000001101;
    16'b0100000010010001: out_v[305] = 10'b0100100111;
    16'b0100100000000000: out_v[305] = 10'b1001101001;
    16'b0100100010010000: out_v[305] = 10'b1001001010;
    16'b0000101010000101: out_v[305] = 10'b0111001001;
    16'b0100100010000000: out_v[305] = 10'b1110001001;
    16'b0110000010000000: out_v[305] = 10'b0001111010;
    16'b0110000010010000: out_v[305] = 10'b1101001010;
    16'b0110000010000001: out_v[305] = 10'b0110011110;
    16'b0100000010010000: out_v[305] = 10'b1100011111;
    16'b0100101010010001: out_v[305] = 10'b1001111110;
    16'b0000101010010001: out_v[305] = 10'b0110011011;
    16'b0100000010000001: out_v[305] = 10'b1011010101;
    16'b0000111010000100: out_v[305] = 10'b1110101001;
    16'b0110000010010001: out_v[305] = 10'b0000111011;
    16'b0110000000000000: out_v[305] = 10'b1101001110;
    16'b0000100010000001: out_v[305] = 10'b1101001010;
    16'b0000000010010001: out_v[305] = 10'b1011010010;
    16'b0100101010000000: out_v[305] = 10'b1111001011;
    16'b0100000000010000: out_v[305] = 10'b0100101111;
    16'b0100101010000001: out_v[305] = 10'b1001100000;
    16'b0000100010010000: out_v[305] = 10'b1001010011;
    16'b0000100000010000: out_v[305] = 10'b1110001011;
    16'b0100101000010000: out_v[305] = 10'b1010100110;
    16'b0100101010010000: out_v[305] = 10'b0111010001;
    16'b0001000010000000: out_v[305] = 10'b0010110101;
    16'b0100100000010000: out_v[305] = 10'b0111011010;
    16'b0010000000010000: out_v[305] = 10'b1100011010;
    16'b0100101000000000: out_v[305] = 10'b1000010110;
    16'b0000000010010000: out_v[305] = 10'b1011001000;
    16'b0000000000001001: out_v[305] = 10'b0100011000;
    16'b0000000000001000: out_v[305] = 10'b1110011010;
    16'b0000001000001000: out_v[305] = 10'b1100110011;
    16'b0001001010000000: out_v[305] = 10'b0110110111;
    16'b0000101000001000: out_v[305] = 10'b1110111010;
    16'b0000001010010000: out_v[305] = 10'b1101110101;
    16'b0100001010010000: out_v[305] = 10'b0100010101;
    16'b0100100000000001: out_v[305] = 10'b0111011010;
    16'b0100101000000001: out_v[305] = 10'b1101011111;
    16'b0000101000001001: out_v[305] = 10'b1010011111;
    16'b0000101010001000: out_v[305] = 10'b0011110010;
    16'b0000001000001001: out_v[305] = 10'b1011100110;
    16'b0000101010001001: out_v[305] = 10'b1101010010;
    16'b0110000000010000: out_v[305] = 10'b0101110011;
    16'b0000100000001001: out_v[305] = 10'b1001100111;
    16'b0011101010010000: out_v[305] = 10'b0001001111;
    16'b0000101001000000: out_v[305] = 10'b1101101011;
    16'b0000001010010001: out_v[305] = 10'b1011010110;
    16'b0000001000010000: out_v[305] = 10'b0111011011;
    16'b0000000000010001: out_v[305] = 10'b0011011010;
    16'b0100001000010000: out_v[305] = 10'b0110111001;
    16'b0000001000010001: out_v[305] = 10'b1101110011;
    16'b0000001010001001: out_v[305] = 10'b0111100001;
    default: out_v[305] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000000000000: out_v[306] = 10'b0100100111;
    16'b0001001000010001: out_v[306] = 10'b1000000111;
    16'b0001000000010001: out_v[306] = 10'b0110000101;
    16'b0000000000010001: out_v[306] = 10'b0100000011;
    16'b0001000000010000: out_v[306] = 10'b0111000101;
    16'b0000001000010001: out_v[306] = 10'b1100010011;
    16'b0000000000000001: out_v[306] = 10'b0110100011;
    16'b0001000000000001: out_v[306] = 10'b1100011110;
    16'b0001000000000000: out_v[306] = 10'b0010011000;
    16'b0000000000010000: out_v[306] = 10'b0100100011;
    16'b0000001000000001: out_v[306] = 10'b1011000011;
    16'b0001001000010000: out_v[306] = 10'b0001110110;
    16'b0001000010010001: out_v[306] = 10'b1101000000;
    16'b0000001010010000: out_v[306] = 10'b1000000110;
    16'b0000000010010000: out_v[306] = 10'b1001100110;
    16'b0000000010000000: out_v[306] = 10'b1100011100;
    16'b0001000010000000: out_v[306] = 10'b0100011010;
    16'b0000001010000000: out_v[306] = 10'b0100110010;
    16'b0001000010010000: out_v[306] = 10'b1100110000;
    16'b0000000010010100: out_v[306] = 10'b1101010010;
    16'b0001000010010100: out_v[306] = 10'b0110000111;
    16'b0001001000000000: out_v[306] = 10'b0010110010;
    16'b0001000000010100: out_v[306] = 10'b1100111100;
    16'b0010000010010000: out_v[306] = 10'b1101111010;
    16'b0000000000010100: out_v[306] = 10'b0000011101;
    16'b0001001010000000: out_v[306] = 10'b0111010000;
    16'b0011000000010000: out_v[306] = 10'b1011011111;
    16'b0011000010010000: out_v[306] = 10'b1001010101;
    16'b0001001000000001: out_v[306] = 10'b0110011001;
    16'b0000001000010000: out_v[306] = 10'b0001111100;
    16'b0001001010010000: out_v[306] = 10'b0000101100;
    16'b0001000010000100: out_v[306] = 10'b1100011111;
    16'b0000000110000000: out_v[306] = 10'b0000011111;
    16'b0001001010010001: out_v[306] = 10'b0111001011;
    16'b0001000010000001: out_v[306] = 10'b1111000110;
    16'b0000001000000000: out_v[306] = 10'b1001111100;
    16'b0000000010010001: out_v[306] = 10'b0001011010;
    16'b0001000000010101: out_v[306] = 10'b1111100010;
    16'b0001000010010101: out_v[306] = 10'b0111100000;
    16'b0000000010010101: out_v[306] = 10'b0011110100;
    16'b0101000010000000: out_v[306] = 10'b1100000000;
    16'b0101000000000000: out_v[306] = 10'b1000001110;
    16'b0000000010000001: out_v[306] = 10'b1111110000;
    16'b0001001010000001: out_v[306] = 10'b0100011010;
    16'b0000001010010001: out_v[306] = 10'b0101011000;
    16'b0000001010000001: out_v[306] = 10'b0000011111;
    default: out_v[306] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010001000000000: out_v[307] = 10'b0000100011;
    16'b0000000000000000: out_v[307] = 10'b0011101000;
    16'b0010011000000000: out_v[307] = 10'b1100110111;
    16'b0010001010000000: out_v[307] = 10'b0100101001;
    16'b1010001000000000: out_v[307] = 10'b0010010100;
    16'b1010010000000000: out_v[307] = 10'b0010010111;
    16'b0000010000000000: out_v[307] = 10'b0010001101;
    16'b0010010000000000: out_v[307] = 10'b0100001001;
    16'b0000001000000000: out_v[307] = 10'b0011110011;
    16'b0010011010000000: out_v[307] = 10'b1001110000;
    16'b0010000000000000: out_v[307] = 10'b0110010011;
    16'b1010001010000000: out_v[307] = 10'b1010001010;
    16'b1010000000000000: out_v[307] = 10'b0101011100;
    16'b1000001000000000: out_v[307] = 10'b0100110010;
    16'b1010011000000000: out_v[307] = 10'b0101000001;
    16'b0000001010000000: out_v[307] = 10'b1111000000;
    16'b0010000010000000: out_v[307] = 10'b1001110010;
    16'b1010001010001000: out_v[307] = 10'b0101000100;
    16'b1010000010001000: out_v[307] = 10'b0101010110;
    16'b1000000000001000: out_v[307] = 10'b0010100011;
    16'b0010000000001000: out_v[307] = 10'b1011111001;
    16'b0010000010001000: out_v[307] = 10'b0111011101;
    16'b1010000000001000: out_v[307] = 10'b0101000010;
    16'b1000000010001000: out_v[307] = 10'b0010011010;
    16'b0010001010001000: out_v[307] = 10'b1110010010;
    16'b1000000000000000: out_v[307] = 10'b1000111000;
    16'b0000000000001000: out_v[307] = 10'b0001101100;
    16'b1011000010001000: out_v[307] = 10'b0101110101;
    16'b1010000010000000: out_v[307] = 10'b1000101101;
    16'b1010001000001000: out_v[307] = 10'b0000100100;
    16'b0010001000001000: out_v[307] = 10'b1100000110;
    16'b1011001010001000: out_v[307] = 10'b0010001100;
    16'b1010000010001010: out_v[307] = 10'b1111000111;
    16'b0000000010001000: out_v[307] = 10'b1001011010;
    16'b1010001010001010: out_v[307] = 10'b1011000101;
    16'b1000001010000000: out_v[307] = 10'b1110000000;
    16'b1000001010001000: out_v[307] = 10'b1000111000;
    16'b1000001000001000: out_v[307] = 10'b0000011000;
    16'b1000000010000000: out_v[307] = 10'b1010110010;
    16'b0000001010001000: out_v[307] = 10'b1101001000;
    16'b0000000010000000: out_v[307] = 10'b1000100111;
    16'b0000000000000010: out_v[307] = 10'b1100011000;
    16'b0000000010000010: out_v[307] = 10'b1111000100;
    16'b0010000010000010: out_v[307] = 10'b1101101000;
    16'b0010001010000010: out_v[307] = 10'b1100101010;
    16'b0010000000000010: out_v[307] = 10'b1000111011;
    16'b0000001010000010: out_v[307] = 10'b1100110110;
    16'b0100001010001000: out_v[307] = 10'b1011000111;
    16'b0000001000001000: out_v[307] = 10'b1100011110;
    16'b0100000010001000: out_v[307] = 10'b0011011001;
    16'b0100000010000000: out_v[307] = 10'b1011010011;
    16'b0100001010000000: out_v[307] = 10'b0110010111;
    16'b0100001000001000: out_v[307] = 10'b0001011111;
    16'b1010011010001000: out_v[307] = 10'b1001110000;
    16'b1010011010000000: out_v[307] = 10'b1000100110;
    16'b0000001010010000: out_v[307] = 10'b1110011101;
    16'b0100001010010000: out_v[307] = 10'b0110100111;
    16'b1100001010001000: out_v[307] = 10'b0011110110;
    default: out_v[307] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001001000000000: out_v[308] = 10'b1101001000;
    16'b0001001000100011: out_v[308] = 10'b1010010111;
    16'b0001001001000011: out_v[308] = 10'b0110000101;
    16'b0001001000000011: out_v[308] = 10'b1010100101;
    16'b0001000000000000: out_v[308] = 10'b1100011111;
    16'b0001000001000011: out_v[308] = 10'b0001110110;
    16'b0001000000000011: out_v[308] = 10'b1001100011;
    16'b0001000001000001: out_v[308] = 10'b0001010111;
    16'b0000000001000000: out_v[308] = 10'b1010000101;
    16'b0000000000000011: out_v[308] = 10'b0101010111;
    16'b0001000001000000: out_v[308] = 10'b0001000111;
    16'b0000000001000011: out_v[308] = 10'b0101011001;
    16'b0001001001100011: out_v[308] = 10'b0111111011;
    16'b0000001000100011: out_v[308] = 10'b0111000101;
    16'b0001001000100000: out_v[308] = 10'b1101001101;
    16'b0001001000010011: out_v[308] = 10'b1111110100;
    16'b0000001000000011: out_v[308] = 10'b1110110001;
    16'b0001001000000001: out_v[308] = 10'b1110111100;
    16'b0001001000100001: out_v[308] = 10'b0000111001;
    16'b0001001010000111: out_v[308] = 10'b1011001101;
    16'b0000000001000001: out_v[308] = 10'b0011111110;
    16'b0001001001000001: out_v[308] = 10'b0010010111;
    16'b0000001001100011: out_v[308] = 10'b0110101100;
    16'b0001000000000001: out_v[308] = 10'b0010001101;
    16'b0000000000100011: out_v[308] = 10'b1100001110;
    16'b0000001001000000: out_v[308] = 10'b1100011011;
    16'b0000001001100000: out_v[308] = 10'b1010000011;
    16'b0000000001000010: out_v[308] = 10'b0110010111;
    16'b0001001011000111: out_v[308] = 10'b1011111101;
    16'b0001000000100011: out_v[308] = 10'b1001001111;
    16'b0000001001000001: out_v[308] = 10'b1110011011;
    16'b0001001000000010: out_v[308] = 10'b0101111001;
    16'b0000001001000011: out_v[308] = 10'b0100110111;
    16'b0000000001100011: out_v[308] = 10'b0111001011;
    16'b0000001000000000: out_v[308] = 10'b1001110010;
    16'b0000000000000000: out_v[308] = 10'b0001100110;
    16'b0000000000100000: out_v[308] = 10'b1000100000;
    16'b0001000000100000: out_v[308] = 10'b1101011010;
    16'b0000001000010000: out_v[308] = 10'b0010110110;
    16'b0000001010010000: out_v[308] = 10'b1001110011;
    16'b0000000000010000: out_v[308] = 10'b1000001110;
    16'b0001000000010000: out_v[308] = 10'b1100110101;
    16'b0000000010000100: out_v[308] = 10'b0100111101;
    16'b0000001010000000: out_v[308] = 10'b1101101000;
    16'b0000000010010000: out_v[308] = 10'b0110100100;
    16'b0001001000010000: out_v[308] = 10'b1001101011;
    16'b0001000010010100: out_v[308] = 10'b1000111111;
    16'b0001000010000100: out_v[308] = 10'b0011110101;
    16'b0000000010010100: out_v[308] = 10'b1011100110;
    16'b0001000000010011: out_v[308] = 10'b1011001111;
    16'b0001000000010001: out_v[308] = 10'b0011100100;
    16'b0001000010010000: out_v[308] = 10'b1000011110;
    16'b0000000000000001: out_v[308] = 10'b0110011001;
    16'b0001000010000000: out_v[308] = 10'b0000011111;
    16'b0001001010010000: out_v[308] = 10'b1111001100;
    16'b0000000010000000: out_v[308] = 10'b0101111111;
    16'b0000000000000100: out_v[308] = 10'b0000010111;
    16'b0001001010000000: out_v[308] = 10'b0110011010;
    16'b0001001010000100: out_v[308] = 10'b0110010100;
    16'b0001000000000100: out_v[308] = 10'b1110100111;
    16'b0001000000000010: out_v[308] = 10'b1000111110;
    16'b0000001010100100: out_v[308] = 10'b0001111110;
    16'b0000001010100000: out_v[308] = 10'b1000101001;
    16'b0000001010000100: out_v[308] = 10'b1010100011;
    16'b0000001010000010: out_v[308] = 10'b1111001011;
    16'b0000001000100000: out_v[308] = 10'b0001110010;
    16'b0000001010000110: out_v[308] = 10'b1011111000;
    16'b0001001010100100: out_v[308] = 10'b1001101010;
    16'b0001001010100000: out_v[308] = 10'b0100011001;
    16'b0000001000010010: out_v[308] = 10'b1011011110;
    16'b0000001010010010: out_v[308] = 10'b1010111011;
    16'b0000000000000010: out_v[308] = 10'b1111110000;
    16'b0001000000100001: out_v[308] = 10'b1111110010;
    16'b0000001000000001: out_v[308] = 10'b1100110010;
    16'b0001000010000111: out_v[308] = 10'b0000010111;
    16'b0000001000000010: out_v[308] = 10'b1111100110;
    16'b0001000001000010: out_v[308] = 10'b0100011101;
    16'b0001000000100010: out_v[308] = 10'b0111101011;
    16'b0000001100000000: out_v[308] = 10'b1000100101;
    16'b0000000100000000: out_v[308] = 10'b1011101100;
    16'b0000000000010011: out_v[308] = 10'b1001110110;
    16'b0000000000010010: out_v[308] = 10'b1011001111;
    16'b0001000011010101: out_v[308] = 10'b1111111001;
    16'b0001000001010011: out_v[308] = 10'b0011101110;
    16'b0001000000100101: out_v[308] = 10'b0000100010;
    16'b0001000000100100: out_v[308] = 10'b1011011001;
    16'b0001001000000100: out_v[308] = 10'b0110000010;
    16'b0001001000000101: out_v[308] = 10'b1001011010;
    16'b0001000010100100: out_v[308] = 10'b1011110001;
    16'b0001001010000101: out_v[308] = 10'b1001001010;
    16'b0001000010100000: out_v[308] = 10'b1111001011;
    16'b0001001000000111: out_v[308] = 10'b1000011111;
    16'b0001000010100001: out_v[308] = 10'b1111000011;
    16'b0000001000000100: out_v[308] = 10'b0111111001;
    16'b0001000010100101: out_v[308] = 10'b0110110111;
    16'b0001000000000101: out_v[308] = 10'b0111110000;
    16'b0000000000100001: out_v[308] = 10'b0110011110;
    16'b0000001000100001: out_v[308] = 10'b0100011000;
    default: out_v[308] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100111010001010: out_v[309] = 10'b1011001011;
    16'b0100111010101010: out_v[309] = 10'b1111011100;
    16'b0100101000101010: out_v[309] = 10'b0001000011;
    16'b0100111010110110: out_v[309] = 10'b0001100110;
    16'b0100111000100110: out_v[309] = 10'b1000110000;
    16'b0100111000110010: out_v[309] = 10'b1010101010;
    16'b0100110010011010: out_v[309] = 10'b1011010011;
    16'b0100111010101110: out_v[309] = 10'b1001011001;
    16'b0100111010111110: out_v[309] = 10'b0111010011;
    16'b0100111000100010: out_v[309] = 10'b0010011110;
    16'b0000101000100010: out_v[309] = 10'b1001010001;
    16'b0100101010101010: out_v[309] = 10'b1111101010;
    16'b0100101010100010: out_v[309] = 10'b0101100011;
    16'b0100101010101110: out_v[309] = 10'b0110110011;
    16'b0100111000110110: out_v[309] = 10'b1100110011;
    16'b0100111010110010: out_v[309] = 10'b1110010011;
    16'b0100111010010110: out_v[309] = 10'b0101010111;
    16'b0100111010111010: out_v[309] = 10'b1001000001;
    16'b0100101000100010: out_v[309] = 10'b0011100011;
    16'b0100111010011010: out_v[309] = 10'b1111010101;
    16'b0100111010101000: out_v[309] = 10'b0110011010;
    16'b0100111010011110: out_v[309] = 10'b1011010101;
    16'b0000101010101000: out_v[309] = 10'b1111111010;
    16'b0100111000101010: out_v[309] = 10'b0010001010;
    16'b0000101010101010: out_v[309] = 10'b1000101111;
    16'b0000101100000010: out_v[309] = 10'b0010110011;
    16'b0100111010100010: out_v[309] = 10'b1110001001;
    16'b0100101000110010: out_v[309] = 10'b0010011011;
    16'b0100111010100110: out_v[309] = 10'b1001111011;
    16'b0100101000100110: out_v[309] = 10'b1011011010;
    16'b0100110010011110: out_v[309] = 10'b0011111011;
    16'b0000000000011100: out_v[309] = 10'b0101000011;
    16'b0000010000010000: out_v[309] = 10'b1101100011;
    16'b0000010000000100: out_v[309] = 10'b1101000001;
    16'b0000010000000000: out_v[309] = 10'b0100010011;
    16'b0000000000010100: out_v[309] = 10'b0111110101;
    16'b0000010000010100: out_v[309] = 10'b0000110111;
    16'b0000000010011100: out_v[309] = 10'b1100010010;
    16'b0000010000011100: out_v[309] = 10'b1001010111;
    16'b0000000010011000: out_v[309] = 10'b0011010011;
    16'b0000000010010100: out_v[309] = 10'b0011110101;
    16'b0000000010010000: out_v[309] = 10'b0000011011;
    16'b0000010010011100: out_v[309] = 10'b1000110100;
    16'b0000000000000000: out_v[309] = 10'b1000011010;
    16'b0000010100010100: out_v[309] = 10'b1001111101;
    16'b0000000110010100: out_v[309] = 10'b1110110101;
    16'b0000000100010100: out_v[309] = 10'b0010110111;
    16'b0000000010011110: out_v[309] = 10'b1010010111;
    16'b0000000010000100: out_v[309] = 10'b1010010010;
    16'b0000000110011100: out_v[309] = 10'b0111001110;
    16'b0000010100110100: out_v[309] = 10'b1000011101;
    16'b0000000010001110: out_v[309] = 10'b1010001100;
    16'b0000000010001100: out_v[309] = 10'b0011110010;
    16'b0000000100010110: out_v[309] = 10'b1101101000;
    16'b0000000000010110: out_v[309] = 10'b1011100001;
    16'b0000010010101110: out_v[309] = 10'b0011011111;
    16'b0000000000001110: out_v[309] = 10'b0011100100;
    16'b0000100010001110: out_v[309] = 10'b1001101111;
    16'b0000000000010000: out_v[309] = 10'b1000011101;
    16'b0000000010000110: out_v[309] = 10'b0011111011;
    16'b0000000010010110: out_v[309] = 10'b1101000101;
    16'b0000000110001110: out_v[309] = 10'b1001000110;
    16'b0000010110010100: out_v[309] = 10'b1000011101;
    16'b0000000110010110: out_v[309] = 10'b0000111000;
    16'b0000000100000100: out_v[309] = 10'b1000110111;
    16'b0000000110000110: out_v[309] = 10'b0111101111;
    16'b0000000010101100: out_v[309] = 10'b0001111111;
    16'b0000000110001100: out_v[309] = 10'b1011001110;
    16'b0000010000010110: out_v[309] = 10'b1100110001;
    16'b0000010010011110: out_v[309] = 10'b1101110111;
    16'b0000000010000010: out_v[309] = 10'b1010010100;
    16'b0000010100010110: out_v[309] = 10'b1101101000;
    16'b0000000110000100: out_v[309] = 10'b1111001100;
    16'b0000010010001110: out_v[309] = 10'b1001111000;
    16'b0000101010001110: out_v[309] = 10'b1101100110;
    16'b0000000010101110: out_v[309] = 10'b0011011111;
    16'b0000000110010000: out_v[309] = 10'b1011010011;
    16'b0100000010010000: out_v[309] = 10'b1011101000;
    16'b0000010100000000: out_v[309] = 10'b1100011100;
    16'b0100010110010000: out_v[309] = 10'b0111111111;
    16'b0100010100010000: out_v[309] = 10'b0101011011;
    16'b0100010010010000: out_v[309] = 10'b0001100110;
    16'b0000000110001000: out_v[309] = 10'b1010001001;
    16'b0000010100010000: out_v[309] = 10'b0001110011;
    16'b0100101010010000: out_v[309] = 10'b0101011111;
    16'b0100010000010000: out_v[309] = 10'b1010101001;
    16'b0000010010011000: out_v[309] = 10'b0111000001;
    16'b0100000100010000: out_v[309] = 10'b0001011111;
    16'b0000000100010000: out_v[309] = 10'b0010101011;
    16'b0000000100000000: out_v[309] = 10'b0011101010;
    16'b0000010010010000: out_v[309] = 10'b1110010000;
    16'b0100010010011000: out_v[309] = 10'b1010100110;
    16'b0100101110010000: out_v[309] = 10'b0011010111;
    16'b0100101100010000: out_v[309] = 10'b1001011111;
    16'b0000000010001000: out_v[309] = 10'b1001111011;
    16'b0100101010011000: out_v[309] = 10'b1001011110;
    16'b0000000000011000: out_v[309] = 10'b1111010111;
    16'b0000000100011000: out_v[309] = 10'b1011011111;
    16'b0000000110000000: out_v[309] = 10'b1000111001;
    16'b0100000010011000: out_v[309] = 10'b1011011111;
    16'b0100000010011100: out_v[309] = 10'b0110001010;
    16'b0000000110011000: out_v[309] = 10'b1110110111;
    16'b0100000000010000: out_v[309] = 10'b0000011101;
    16'b0100010100000000: out_v[309] = 10'b0001001101;
    16'b0000010100110000: out_v[309] = 10'b0001011010;
    16'b0100000110010000: out_v[309] = 10'b1111110110;
    16'b0100111100010000: out_v[309] = 10'b1010010000;
    16'b0000010110010000: out_v[309] = 10'b0111110011;
    16'b0100000110011000: out_v[309] = 10'b0011110111;
    16'b0100101110011000: out_v[309] = 10'b0011101111;
    16'b0100010000000000: out_v[309] = 10'b1100001101;
    16'b0100101000100000: out_v[309] = 10'b0000110101;
    16'b0100101100110010: out_v[309] = 10'b0001111101;
    16'b0100101000111110: out_v[309] = 10'b0010010001;
    16'b0000101100010010: out_v[309] = 10'b1001000100;
    16'b0100101000110110: out_v[309] = 10'b1001001011;
    16'b0000101100100010: out_v[309] = 10'b0111111110;
    16'b0100000000110100: out_v[309] = 10'b0101010100;
    16'b0100101000100100: out_v[309] = 10'b0000110011;
    16'b0100101100100010: out_v[309] = 10'b0110111110;
    16'b0000101000010010: out_v[309] = 10'b0010010101;
    16'b0100111000000110: out_v[309] = 10'b0001010110;
    16'b0000101100001010: out_v[309] = 10'b0111000010;
    16'b0100101000110000: out_v[309] = 10'b0001001111;
    16'b0100101000101110: out_v[309] = 10'b0011001001;
    16'b0100101000111000: out_v[309] = 10'b1011101110;
    16'b0100111000010010: out_v[309] = 10'b1000110111;
    16'b0000101000000010: out_v[309] = 10'b1000110011;
    16'b0100111000100100: out_v[309] = 10'b0100111111;
    16'b0000101100011010: out_v[309] = 10'b1111001000;
    16'b0100000000110000: out_v[309] = 10'b1101010001;
    16'b0100110000010010: out_v[309] = 10'b0101110110;
    16'b0100101000111010: out_v[309] = 10'b1011000011;
    16'b0100000000100000: out_v[309] = 10'b1001110110;
    16'b0000101000101010: out_v[309] = 10'b1011100010;
    16'b0100101100110000: out_v[309] = 10'b0010110110;
    16'b0000101000100110: out_v[309] = 10'b1100111011;
    16'b0100101000101000: out_v[309] = 10'b0101011110;
    16'b0100010010101000: out_v[309] = 10'b1011110010;
    16'b0100000000101000: out_v[309] = 10'b0010110111;
    16'b0100010010010100: out_v[309] = 10'b0101111000;
    16'b0100101010101000: out_v[309] = 10'b0011101001;
    16'b0100111000100000: out_v[309] = 10'b0000110110;
    16'b0100000100100000: out_v[309] = 10'b1011100011;
    16'b0100111010110000: out_v[309] = 10'b1000100110;
    16'b0100111010100000: out_v[309] = 10'b0011011110;
    16'b0100010000101000: out_v[309] = 10'b1010100110;
    16'b0100010010100000: out_v[309] = 10'b0001111110;
    16'b0100010000100000: out_v[309] = 10'b1110000101;
    16'b0100111010110100: out_v[309] = 10'b0011011010;
    16'b0100010000010100: out_v[309] = 10'b1010101111;
    16'b0100111000101000: out_v[309] = 10'b1011011110;
    16'b0100010010110100: out_v[309] = 10'b0101111011;
    16'b0100010010110000: out_v[309] = 10'b1111001000;
    16'b0100001010101000: out_v[309] = 10'b1110011011;
    16'b0100000010101000: out_v[309] = 10'b1111000010;
    16'b0100111000110000: out_v[309] = 10'b1011100101;
    16'b0100010010111000: out_v[309] = 10'b0011111011;
    16'b0000010010010100: out_v[309] = 10'b1110011001;
    16'b0000010010001000: out_v[309] = 10'b0110110011;
    16'b0100010010001000: out_v[309] = 10'b1101110111;
    16'b0100111000101110: out_v[309] = 10'b1011001110;
    16'b0100010000000110: out_v[309] = 10'b1001101001;
    16'b0000010000001000: out_v[309] = 10'b0000110101;
    16'b1000101100000110: out_v[309] = 10'b0111000011;
    16'b0100010000100110: out_v[309] = 10'b0010111110;
    16'b0100101100100110: out_v[309] = 10'b0111001110;
    16'b0000010000011110: out_v[309] = 10'b1000101110;
    16'b0100010000100100: out_v[309] = 10'b0001111101;
    16'b0100010000000100: out_v[309] = 10'b1000110100;
    16'b0100000000100100: out_v[309] = 10'b1001001011;
    16'b0100010000001110: out_v[309] = 10'b1101111011;
    16'b0100010000001100: out_v[309] = 10'b1011101010;
    16'b1100101000100110: out_v[309] = 10'b1011111001;
    16'b0000101100000110: out_v[309] = 10'b1001011001;
    16'b0100000000000100: out_v[309] = 10'b1001001000;
    16'b0100000000100110: out_v[309] = 10'b1110111110;
    16'b0000010000001100: out_v[309] = 10'b0101011001;
    16'b0100111000001110: out_v[309] = 10'b1000101110;
    16'b1100101100100110: out_v[309] = 10'b0001010101;
    16'b0100110000100110: out_v[309] = 10'b1111110101;
    16'b0100110000011110: out_v[309] = 10'b0111100010;
    16'b0100010000011110: out_v[309] = 10'b0011010111;
    16'b0000000000000100: out_v[309] = 10'b0111101001;
    16'b0000101100100110: out_v[309] = 10'b0110111111;
    16'b0000101100010110: out_v[309] = 10'b0111010010;
    16'b0100100000100110: out_v[309] = 10'b1101110011;
    16'b0100101100110110: out_v[309] = 10'b0001011010;
    16'b0100110000000110: out_v[309] = 10'b1101111110;
    16'b0100110000001110: out_v[309] = 10'b1110101111;
    16'b0100011000110100: out_v[309] = 10'b0101000111;
    16'b0000010000110000: out_v[309] = 10'b0101011010;
    16'b0000010000100100: out_v[309] = 10'b0110110010;
    16'b0000010000110100: out_v[309] = 10'b0110101001;
    16'b0100011000110000: out_v[309] = 10'b1101100111;
    16'b0100111000110100: out_v[309] = 10'b0110000110;
    16'b0100010000110100: out_v[309] = 10'b0010100110;
    16'b0100010000110000: out_v[309] = 10'b1111100001;
    16'b0100010100110000: out_v[309] = 10'b1001110100;
    16'b0100011000100100: out_v[309] = 10'b0111011011;
    16'b0000010000100000: out_v[309] = 10'b0011011110;
    16'b0000010100100100: out_v[309] = 10'b0010011011;
    16'b0000111000110000: out_v[309] = 10'b1101001110;
    16'b0000010100000100: out_v[309] = 10'b1000100101;
    16'b0100111100110010: out_v[309] = 10'b0011101011;
    16'b0100010100110100: out_v[309] = 10'b1110000001;
    16'b0000000000110000: out_v[309] = 10'b0110011001;
    16'b0100111100110000: out_v[309] = 10'b0011100111;
    16'b0000011000110000: out_v[309] = 10'b0111100111;
    16'b0000010010011010: out_v[309] = 10'b1111100000;
    16'b0100010000111100: out_v[309] = 10'b0111000001;
    16'b0100000000111100: out_v[309] = 10'b1100010011;
    16'b0000010010001100: out_v[309] = 10'b1110110001;
    16'b0100000010101100: out_v[309] = 10'b1111000101;
    16'b0100000100110100: out_v[309] = 10'b1101010111;
    16'b0000000000110100: out_v[309] = 10'b0101110100;
    16'b0100000000111000: out_v[309] = 10'b1100000011;
    16'b0100000010111000: out_v[309] = 10'b1100100011;
    16'b0000000000100100: out_v[309] = 10'b0110001010;
    16'b0100000100100100: out_v[309] = 10'b0110001011;
    16'b0100010010101100: out_v[309] = 10'b1111100000;
    16'b0100000000101100: out_v[309] = 10'b0111001011;
    16'b0100010000101100: out_v[309] = 10'b0011100101;
    16'b0100001000110000: out_v[309] = 10'b1001000011;
    16'b0000111000110010: out_v[309] = 10'b1000100010;
    16'b0000111000100000: out_v[309] = 10'b1101101111;
    16'b0000111100010010: out_v[309] = 10'b1000010111;
    16'b0000101000110000: out_v[309] = 10'b1101000111;
    16'b0000101000110010: out_v[309] = 10'b1101010111;
    16'b0000101000100000: out_v[309] = 10'b1001000111;
    16'b0000111000100010: out_v[309] = 10'b1100100100;
    16'b0000111100010000: out_v[309] = 10'b1111000111;
    default: out_v[309] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000111000101: out_v[310] = 10'b0011011001;
    16'b0000000101100001: out_v[310] = 10'b1101110100;
    16'b0000100101100101: out_v[310] = 10'b0001110111;
    16'b0000010101000101: out_v[310] = 10'b1111000010;
    16'b0000000100100001: out_v[310] = 10'b0111111000;
    16'b0000000100100101: out_v[310] = 10'b0111111011;
    16'b0000000100000001: out_v[310] = 10'b0000001110;
    16'b0000000000000001: out_v[310] = 10'b1100111011;
    16'b0000010101100100: out_v[310] = 10'b0110100111;
    16'b0000010101000001: out_v[310] = 10'b1111110011;
    16'b0000000000100001: out_v[310] = 10'b1001000011;
    16'b0000010101100101: out_v[310] = 10'b0000011011;
    16'b0000100100000001: out_v[310] = 10'b1101011110;
    16'b0000000101000101: out_v[310] = 10'b1101001110;
    16'b0000000101100101: out_v[310] = 10'b1110010110;
    16'b0000010100000001: out_v[310] = 10'b0000110111;
    16'b0000010100000101: out_v[310] = 10'b1110010111;
    16'b0000010111100101: out_v[310] = 10'b1101011111;
    16'b0000100100000000: out_v[310] = 10'b0100010101;
    16'b0000010111000101: out_v[310] = 10'b1011000110;
    16'b0000010101100001: out_v[310] = 10'b1011011111;
    16'b0000000111101101: out_v[310] = 10'b0000111101;
    16'b0000000111100101: out_v[310] = 10'b0000011101;
    16'b0000100100100001: out_v[310] = 10'b0111001110;
    16'b0000000101000001: out_v[310] = 10'b1001011111;
    16'b0000010011000101: out_v[310] = 10'b1100111110;
    16'b0000010001000101: out_v[310] = 10'b1110000011;
    16'b0000000100000000: out_v[310] = 10'b0011100110;
    16'b0000000111001101: out_v[310] = 10'b1001101001;
    16'b0000100101000100: out_v[310] = 10'b0100011111;
    16'b0000000101100100: out_v[310] = 10'b1101001011;
    16'b0000000001000101: out_v[310] = 10'b0100000001;
    16'b0000000111100100: out_v[310] = 10'b1011001101;
    16'b0000000100000101: out_v[310] = 10'b1100010010;
    16'b0000010100100001: out_v[310] = 10'b1101010001;
    16'b0000100101000101: out_v[310] = 10'b1100010101;
    16'b0000110101000101: out_v[310] = 10'b1101111110;
    16'b0000000101000100: out_v[310] = 10'b0010101000;
    16'b0000000100100000: out_v[310] = 10'b1000001111;
    16'b0000000000100000: out_v[310] = 10'b1101011001;
    16'b0000000101000000: out_v[310] = 10'b1100100111;
    16'b0000000100000100: out_v[310] = 10'b1001101010;
    16'b0000010100000100: out_v[310] = 10'b0011010100;
    16'b0000000000000000: out_v[310] = 10'b1011000100;
    16'b0000000001000000: out_v[310] = 10'b1010110010;
    16'b0000000101100000: out_v[310] = 10'b1011001000;
    16'b0000010101000000: out_v[310] = 10'b0111110100;
    16'b0000010101100000: out_v[310] = 10'b0010011011;
    16'b0000000000000100: out_v[310] = 10'b1011010011;
    16'b0000000001100000: out_v[310] = 10'b0110010101;
    16'b0000000110000100: out_v[310] = 10'b0110101011;
    16'b0000010100000000: out_v[310] = 10'b0011100010;
    16'b0000010001100000: out_v[310] = 10'b1001101111;
    16'b0000010100100000: out_v[310] = 10'b1110100110;
    16'b0000010000100000: out_v[310] = 10'b1000001100;
    16'b0000001000100001: out_v[310] = 10'b1111011001;
    16'b0000010001000000: out_v[310] = 10'b1011001001;
    16'b0000010000000000: out_v[310] = 10'b0011001100;
    16'b0000010101000100: out_v[310] = 10'b0011010010;
    16'b0000000010000100: out_v[310] = 10'b1001010011;
    16'b0000000100100100: out_v[310] = 10'b0110110101;
    16'b0000010100100100: out_v[310] = 10'b0100110010;
    16'b0000000111101100: out_v[310] = 10'b1001101110;
    16'b0000000100001000: out_v[310] = 10'b0100111110;
    16'b0000010000000001: out_v[310] = 10'b0000000101;
    16'b1000000100101000: out_v[310] = 10'b1101000111;
    16'b0000010000001001: out_v[310] = 10'b1001110011;
    16'b0000010100100101: out_v[310] = 10'b1000110101;
    16'b1000010000100000: out_v[310] = 10'b1110101100;
    16'b1000000100100000: out_v[310] = 10'b1010010111;
    16'b0000000101101100: out_v[310] = 10'b1010110110;
    16'b0000010110100100: out_v[310] = 10'b1011000101;
    16'b0000000100101000: out_v[310] = 10'b1000000110;
    16'b0000010000100001: out_v[310] = 10'b0101001001;
    16'b0000010000100100: out_v[310] = 10'b1100101110;
    16'b0000010000100101: out_v[310] = 10'b1110001101;
    16'b0000000100101001: out_v[310] = 10'b1110100110;
    16'b0000010000000101: out_v[310] = 10'b1010001110;
    16'b0000000111000100: out_v[310] = 10'b0001110100;
    16'b0000000101001100: out_v[310] = 10'b1111100111;
    16'b0000000011101100: out_v[310] = 10'b1100010101;
    16'b0000000110101100: out_v[310] = 10'b0110000000;
    16'b0000000001100100: out_v[310] = 10'b0100101011;
    16'b0000000111001100: out_v[310] = 10'b0011110010;
    16'b0000000101101101: out_v[310] = 10'b0110000011;
    16'b0000000001000100: out_v[310] = 10'b0110001001;
    16'b0000010001100101: out_v[310] = 10'b1110101001;
    16'b0000010001100100: out_v[310] = 10'b1101001000;
    16'b0000010001000100: out_v[310] = 10'b0011100111;
    16'b0000000010100100: out_v[310] = 10'b0101010000;
    16'b0000000001000001: out_v[310] = 10'b1111111010;
    16'b0000000010100000: out_v[310] = 10'b0110010010;
    16'b0000001000000001: out_v[310] = 10'b1000011001;
    16'b0000000010100001: out_v[310] = 10'b0011111110;
    16'b0000000001100001: out_v[310] = 10'b1011000100;
    16'b0000000000100100: out_v[310] = 10'b0111011010;
    16'b0000000000100101: out_v[310] = 10'b0111100010;
    16'b0000001001000001: out_v[310] = 10'b0011101111;
    16'b0000000110100100: out_v[310] = 10'b1011100111;
    16'b0000000001100101: out_v[310] = 10'b1101100011;
    16'b0000000010101001: out_v[310] = 10'b0010111101;
    16'b0000000010101100: out_v[310] = 10'b0100111111;
    16'b0000000000000101: out_v[310] = 10'b1100010011;
    16'b0000000010101101: out_v[310] = 10'b1100100111;
    16'b0000001100000001: out_v[310] = 10'b0011010011;
    16'b0000000010000101: out_v[310] = 10'b0111111010;
    16'b0000000010000001: out_v[310] = 10'b1100110011;
    16'b0000000010100101: out_v[310] = 10'b0011111110;
    16'b0000000000001001: out_v[310] = 10'b0010010010;
    16'b0000000010101000: out_v[310] = 10'b1001110010;
    16'b0000000010001101: out_v[310] = 10'b1010111101;
    16'b0000000010001001: out_v[310] = 10'b0010110001;
    16'b0000001101000001: out_v[310] = 10'b0111010110;
    16'b0000000000101000: out_v[310] = 10'b0001010111;
    16'b0000001111000100: out_v[310] = 10'b1011110001;
    16'b0000100000100001: out_v[310] = 10'b1001100010;
    16'b0000001100000100: out_v[310] = 10'b0110111001;
    16'b0000001101000100: out_v[310] = 10'b1001010110;
    16'b0000001100000000: out_v[310] = 10'b0100001010;
    16'b0000001101100101: out_v[310] = 10'b0101011111;
    16'b0000001101000000: out_v[310] = 10'b1111010110;
    16'b0000001101000101: out_v[310] = 10'b1101101001;
    16'b0000001000000000: out_v[310] = 10'b0010100111;
    16'b0000000110000000: out_v[310] = 10'b0000110110;
    16'b0000010000000100: out_v[310] = 10'b1000110101;
    16'b0000010011000100: out_v[310] = 10'b1011110111;
    16'b0000001001100001: out_v[310] = 10'b1011100101;
    16'b0000010111000100: out_v[310] = 10'b1011010101;
    16'b0000000000001000: out_v[310] = 10'b0101010100;
    16'b0010000000000000: out_v[310] = 10'b1111001011;
    16'b0000000000101001: out_v[310] = 10'b0001101010;
    16'b0000000101101000: out_v[310] = 10'b1011100001;
    16'b0000000000101100: out_v[310] = 10'b1010111011;
    16'b0000000001101000: out_v[310] = 10'b0100111111;
    16'b0000000001101001: out_v[310] = 10'b1010101011;
    16'b0000000101101001: out_v[310] = 10'b1101101000;
    16'b0000000101001001: out_v[310] = 10'b0010100111;
    16'b0000000100001001: out_v[310] = 10'b1110001001;
    16'b0000000100101100: out_v[310] = 10'b1110010001;
    16'b0000000001101101: out_v[310] = 10'b0011010011;
    16'b0000010011100100: out_v[310] = 10'b1101001010;
    16'b0000001101100001: out_v[310] = 10'b1100010110;
    16'b0000001100100001: out_v[310] = 10'b1100010111;
    16'b0000000011100100: out_v[310] = 10'b1111000011;
    16'b0000000110100000: out_v[310] = 10'b1001101011;
    16'b0000000110100101: out_v[310] = 10'b1000110100;
    16'b0000000110000001: out_v[310] = 10'b1101100110;
    16'b0000000110000101: out_v[310] = 10'b0011010100;
    16'b0000000110100001: out_v[310] = 10'b1100100010;
    default: out_v[310] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000001001000: out_v[311] = 10'b1000100111;
    16'b0010101011000000: out_v[311] = 10'b1010101011;
    16'b1000101011001001: out_v[311] = 10'b1011010011;
    16'b0000100001001000: out_v[311] = 10'b1001101011;
    16'b0010101010010000: out_v[311] = 10'b0101000111;
    16'b0000101011001000: out_v[311] = 10'b0011011100;
    16'b0010101010000000: out_v[311] = 10'b0111000101;
    16'b1000111011001001: out_v[311] = 10'b1010010010;
    16'b0000001011000000: out_v[311] = 10'b0101000101;
    16'b0000101011000000: out_v[311] = 10'b1010100111;
    16'b1000111011000001: out_v[311] = 10'b1000001001;
    16'b1000101011001000: out_v[311] = 10'b1111010011;
    16'b0010001011000000: out_v[311] = 10'b1101110000;
    16'b0000101010000000: out_v[311] = 10'b0110111001;
    16'b0000101011001001: out_v[311] = 10'b1010110111;
    16'b0010000001000000: out_v[311] = 10'b0100110110;
    16'b0000000001000000: out_v[311] = 10'b0111000001;
    16'b0000101011011000: out_v[311] = 10'b1101011110;
    16'b0010101011001000: out_v[311] = 10'b0011001110;
    16'b0000001011001000: out_v[311] = 10'b0101010101;
    16'b0010101010001000: out_v[311] = 10'b0111110110;
    16'b1100111011001001: out_v[311] = 10'b1101001100;
    16'b0010101011010000: out_v[311] = 10'b0000110001;
    16'b1000100001001000: out_v[311] = 10'b1111010011;
    16'b1100111011000001: out_v[311] = 10'b0111011111;
    16'b1100101011001001: out_v[311] = 10'b1110101100;
    16'b0010100010000000: out_v[311] = 10'b0111001110;
    16'b0010101010001001: out_v[311] = 10'b0001111110;
    16'b0000101010001000: out_v[311] = 10'b0101000011;
    16'b0010101011001001: out_v[311] = 10'b0101011000;
    16'b1000000001001000: out_v[311] = 10'b1110110001;
    16'b1000000001001001: out_v[311] = 10'b0011000111;
    16'b1010101011001001: out_v[311] = 10'b1011000111;
    16'b0010101011011000: out_v[311] = 10'b1110011001;
    16'b0010001011001000: out_v[311] = 10'b0111011010;
    16'b0000100001000000: out_v[311] = 10'b1111001101;
    16'b0010101000000000: out_v[311] = 10'b1000100101;
    16'b0010100000000000: out_v[311] = 10'b1111100110;
    16'b0010000000000000: out_v[311] = 10'b1111100001;
    16'b1010000000000000: out_v[311] = 10'b0110011101;
    16'b0010001000000000: out_v[311] = 10'b0010110101;
    16'b1000000000000000: out_v[311] = 10'b1011001010;
    16'b0010001001000000: out_v[311] = 10'b0001011010;
    16'b0000101000000000: out_v[311] = 10'b1101010011;
    16'b0000000000000000: out_v[311] = 10'b0001010111;
    16'b1110010000000000: out_v[311] = 10'b1101000100;
    16'b1000001011000000: out_v[311] = 10'b1011011111;
    16'b1100001011000000: out_v[311] = 10'b1011010110;
    16'b1000000001000000: out_v[311] = 10'b0110101001;
    16'b0010010000001001: out_v[311] = 10'b0010110101;
    16'b1010000001000000: out_v[311] = 10'b1010011000;
    16'b1110000000000000: out_v[311] = 10'b0110100110;
    16'b1000111011000000: out_v[311] = 10'b1000010101;
    16'b0000100011000000: out_v[311] = 10'b1010100111;
    16'b1100100011000000: out_v[311] = 10'b1111100111;
    16'b1000000011000000: out_v[311] = 10'b0010110111;
    16'b1010000011000000: out_v[311] = 10'b1010011010;
    16'b1000100011000000: out_v[311] = 10'b1110110110;
    16'b1010001011000000: out_v[311] = 10'b0101001011;
    16'b1000011011000000: out_v[311] = 10'b1110000100;
    16'b1000101011000000: out_v[311] = 10'b0011111110;
    16'b0010000000001000: out_v[311] = 10'b1100000101;
    16'b1010010000000000: out_v[311] = 10'b1110001001;
    16'b1100101011000000: out_v[311] = 10'b1011110101;
    16'b1000011011000001: out_v[311] = 10'b1001001110;
    16'b1100111011000000: out_v[311] = 10'b0111011100;
    16'b0000000011000000: out_v[311] = 10'b1001000100;
    16'b1100011011000000: out_v[311] = 10'b1111110010;
    16'b1110000001000000: out_v[311] = 10'b1010001101;
    16'b0100101011000000: out_v[311] = 10'b0100110100;
    16'b0010010000000001: out_v[311] = 10'b1101100110;
    16'b1010000010000000: out_v[311] = 10'b0010011111;
    16'b0000100010000000: out_v[311] = 10'b1000111110;
    16'b0010000011000000: out_v[311] = 10'b1101110010;
    16'b1010010000000001: out_v[311] = 10'b1100111101;
    16'b1010011001000001: out_v[311] = 10'b0010111001;
    16'b1010001001000000: out_v[311] = 10'b1010001101;
    16'b1010011010000000: out_v[311] = 10'b0011011010;
    16'b1010010001000001: out_v[311] = 10'b1011010111;
    16'b0010101001000000: out_v[311] = 10'b0100010100;
    16'b1000101001000000: out_v[311] = 10'b1011000110;
    16'b1010011001000000: out_v[311] = 10'b1101011011;
    16'b1010111011000000: out_v[311] = 10'b0001011110;
    16'b1010101011000000: out_v[311] = 10'b1111001010;
    16'b1110011000000000: out_v[311] = 10'b1110100100;
    16'b0000101001000000: out_v[311] = 10'b0011010101;
    16'b1010011000000000: out_v[311] = 10'b1110010111;
    16'b1110011011000000: out_v[311] = 10'b1110011001;
    16'b0110010000000001: out_v[311] = 10'b1000001001;
    16'b1110010000000001: out_v[311] = 10'b1001011111;
    16'b1010001000000000: out_v[311] = 10'b0001011001;
    16'b1010011011000000: out_v[311] = 10'b1111011000;
    16'b1010101001000000: out_v[311] = 10'b0011011011;
    16'b1010111001000000: out_v[311] = 10'b0100111000;
    16'b1010010001000000: out_v[311] = 10'b1111111110;
    16'b1110011011000001: out_v[311] = 10'b0111100010;
    16'b1010111011000001: out_v[311] = 10'b1111001010;
    16'b1010001010000000: out_v[311] = 10'b0001110101;
    16'b1010011011000001: out_v[311] = 10'b0011101010;
    16'b0010010000000000: out_v[311] = 10'b0011011001;
    16'b1110010001000000: out_v[311] = 10'b0101111011;
    16'b0000000000001001: out_v[311] = 10'b0100001100;
    16'b0000100000010000: out_v[311] = 10'b1000101111;
    16'b0000100000001000: out_v[311] = 10'b0101110110;
    16'b1000000000001000: out_v[311] = 10'b0101010011;
    16'b0000000000001000: out_v[311] = 10'b1100000111;
    16'b0100110000000001: out_v[311] = 10'b0000111110;
    16'b0000100000000000: out_v[311] = 10'b0001110011;
    16'b0000110000001001: out_v[311] = 10'b1110001011;
    16'b1000000000001001: out_v[311] = 10'b0111111001;
    16'b0000010000000001: out_v[311] = 10'b0101100011;
    16'b0000000000010000: out_v[311] = 10'b1001110011;
    16'b0000010000000000: out_v[311] = 10'b1101001000;
    16'b1000100000001000: out_v[311] = 10'b0000010110;
    16'b0000100000001001: out_v[311] = 10'b0001111010;
    16'b1000100000001001: out_v[311] = 10'b0011101110;
    16'b0000110000000001: out_v[311] = 10'b0011011101;
    16'b0000001000010000: out_v[311] = 10'b0101011011;
    16'b0000010000001001: out_v[311] = 10'b0110110011;
    16'b0100010000000000: out_v[311] = 10'b1000110110;
    16'b0000110000000000: out_v[311] = 10'b0001110011;
    16'b0100110000000000: out_v[311] = 10'b0111010010;
    16'b0000100000000001: out_v[311] = 10'b0101111101;
    16'b0010000001001000: out_v[311] = 10'b1110010010;
    16'b0010000000001001: out_v[311] = 10'b0001100001;
    16'b0100010000000001: out_v[311] = 10'b1100101010;
    16'b0000100000011000: out_v[311] = 10'b0011100110;
    16'b0100000000000000: out_v[311] = 10'b0010010010;
    16'b0100100000000000: out_v[311] = 10'b0101011101;
    16'b0000000000011000: out_v[311] = 10'b0001011010;
    16'b1000110000001001: out_v[311] = 10'b1000111111;
    16'b0010001010000000: out_v[311] = 10'b1111001001;
    16'b0000101010010000: out_v[311] = 10'b1110101010;
    16'b0010000010000000: out_v[311] = 10'b0101100001;
    16'b0010101000010000: out_v[311] = 10'b1001100100;
    16'b0000101000001000: out_v[311] = 10'b0001111011;
    16'b0000101010011000: out_v[311] = 10'b1110010111;
    16'b0000101000010000: out_v[311] = 10'b0011000011;
    16'b0010100010010000: out_v[311] = 10'b1010100101;
    16'b0010101010011000: out_v[311] = 10'b1001110111;
    16'b0010100000010000: out_v[311] = 10'b1101100111;
    16'b0000100010010000: out_v[311] = 10'b0100001111;
    16'b0000101001001000: out_v[311] = 10'b1010111011;
    16'b1000001011001000: out_v[311] = 10'b0000100011;
    16'b0000001001000000: out_v[311] = 10'b1110100100;
    16'b1000010000000001: out_v[311] = 10'b1011000010;
    16'b1000010000001001: out_v[311] = 10'b0011011001;
    16'b0000000011001000: out_v[311] = 10'b0101111000;
    16'b1000000010001001: out_v[311] = 10'b0111101010;
    16'b1010000000001001: out_v[311] = 10'b1101010010;
    16'b1010000000001000: out_v[311] = 10'b1101100010;
    16'b1000000010001000: out_v[311] = 10'b1001000000;
    16'b0010010000101001: out_v[311] = 10'b1010110000;
    16'b0010100000001000: out_v[311] = 10'b1001001000;
    16'b0010100000001001: out_v[311] = 10'b0011011010;
    16'b0010110000001001: out_v[311] = 10'b0001101101;
    16'b0010111000001001: out_v[311] = 10'b0111000110;
    16'b0010000000101000: out_v[311] = 10'b1111110111;
    16'b0000101000001001: out_v[311] = 10'b0101011111;
    16'b0010000000101001: out_v[311] = 10'b1100001111;
    16'b0010101000001000: out_v[311] = 10'b1110110011;
    16'b0010000000000001: out_v[311] = 10'b1001000101;
    16'b0010101000001001: out_v[311] = 10'b0101011111;
    16'b0010100001000000: out_v[311] = 10'b0111011101;
    16'b1010000001001000: out_v[311] = 10'b0101110100;
    16'b0000100001001001: out_v[311] = 10'b1110000110;
    16'b1000100001001001: out_v[311] = 10'b0111001011;
    16'b0010100001001000: out_v[311] = 10'b0010110100;
    16'b0000101011010000: out_v[311] = 10'b1011011011;
    16'b1010000001001001: out_v[311] = 10'b1101110010;
    16'b0110000000001001: out_v[311] = 10'b1011001001;
    16'b0000000000000001: out_v[311] = 10'b1001100111;
    16'b0110000000001000: out_v[311] = 10'b1011001011;
    16'b0100000000001001: out_v[311] = 10'b1101100010;
    16'b0110010000001001: out_v[311] = 10'b0010101100;
    default: out_v[311] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100010000101101: out_v[312] = 10'b0011110110;
    16'b1100010000101100: out_v[312] = 10'b1000010011;
    16'b1100010101101101: out_v[312] = 10'b0100110011;
    16'b1100010000101101: out_v[312] = 10'b0100011111;
    16'b0100010000101100: out_v[312] = 10'b1011001111;
    16'b1010000100001101: out_v[312] = 10'b0110110101;
    16'b1100010000001100: out_v[312] = 10'b0110110011;
    16'b1100010100000101: out_v[312] = 10'b0100110011;
    16'b1100010100001101: out_v[312] = 10'b1100010100;
    16'b1100010000100100: out_v[312] = 10'b1111000010;
    16'b1100010000001101: out_v[312] = 10'b0111111010;
    16'b1000000101001101: out_v[312] = 10'b0111110110;
    16'b1100010000100101: out_v[312] = 10'b0000100010;
    16'b1100010100101100: out_v[312] = 10'b0110010001;
    16'b0100010001101100: out_v[312] = 10'b1011101001;
    16'b1100010100101101: out_v[312] = 10'b1000110011;
    16'b1000010100001101: out_v[312] = 10'b1111110111;
    16'b1110000101001101: out_v[312] = 10'b1100011010;
    16'b1100000101001101: out_v[312] = 10'b0110101011;
    16'b1100000000001100: out_v[312] = 10'b1100100001;
    16'b1010000101001101: out_v[312] = 10'b1110000011;
    16'b0010000100001101: out_v[312] = 10'b1001011111;
    16'b1100000000001101: out_v[312] = 10'b0100000011;
    16'b0100000000101100: out_v[312] = 10'b1110111011;
    16'b1000010101001101: out_v[312] = 10'b1111111000;
    16'b0100010000101000: out_v[312] = 10'b1010001111;
    16'b1100010001101101: out_v[312] = 10'b0011001010;
    16'b0100010001101101: out_v[312] = 10'b0100010011;
    16'b1100000100001101: out_v[312] = 10'b1101000111;
    16'b1100010000101000: out_v[312] = 10'b1111000011;
    16'b1000000100001101: out_v[312] = 10'b1001000001;
    16'b1000000101001001: out_v[312] = 10'b1010110001;
    16'b0100010000100100: out_v[312] = 10'b1110100110;
    16'b1110000100001101: out_v[312] = 10'b0110011011;
    16'b0100000000101000: out_v[312] = 10'b1100001001;
    16'b1100010000100000: out_v[312] = 10'b1111000010;
    16'b1100010101001101: out_v[312] = 10'b1101101111;
    16'b0100000000100000: out_v[312] = 10'b0010110001;
    16'b1100010001001101: out_v[312] = 10'b1001100010;
    16'b1000010100101101: out_v[312] = 10'b1011101011;
    16'b1100000001001101: out_v[312] = 10'b1110111011;
    16'b1100000100000101: out_v[312] = 10'b0101100000;
    16'b1010000101001001: out_v[312] = 10'b1100001011;
    16'b1100010100100101: out_v[312] = 10'b1100001100;
    16'b1000000100001001: out_v[312] = 10'b0010010111;
    16'b0000000000001000: out_v[312] = 10'b1100100111;
    16'b0000000000000000: out_v[312] = 10'b0001101011;
    16'b0000000001000000: out_v[312] = 10'b0010001101;
    16'b0000000001000100: out_v[312] = 10'b1010100010;
    16'b0000000000000100: out_v[312] = 10'b1110101101;
    16'b0000000000000101: out_v[312] = 10'b0010011100;
    16'b0100000000000100: out_v[312] = 10'b0001110010;
    16'b0000000001000101: out_v[312] = 10'b1001010111;
    16'b0000010001000000: out_v[312] = 10'b1000000110;
    16'b1000010001101000: out_v[312] = 10'b1000000110;
    16'b0000010001100001: out_v[312] = 10'b0011111111;
    16'b0000010001101000: out_v[312] = 10'b1111010010;
    16'b0000010001001000: out_v[312] = 10'b1001100101;
    16'b0000000000101101: out_v[312] = 10'b1011011011;
    16'b0000000001101101: out_v[312] = 10'b1111110110;
    16'b0000000001001000: out_v[312] = 10'b0000110110;
    16'b0000000001101000: out_v[312] = 10'b1011100110;
    16'b0000010001100000: out_v[312] = 10'b1110000101;
    16'b1000000000101000: out_v[312] = 10'b0000001100;
    16'b0000000000101000: out_v[312] = 10'b1110000111;
    16'b0000010001101001: out_v[312] = 10'b1111001011;
    16'b0000010001101101: out_v[312] = 10'b0100110010;
    16'b1000010000100101: out_v[312] = 10'b1100000010;
    16'b1000000001100000: out_v[312] = 10'b1000101011;
    16'b0000000000101100: out_v[312] = 10'b0010101110;
    16'b1000010001101101: out_v[312] = 10'b1110110110;
    16'b0000010000101100: out_v[312] = 10'b1010001110;
    16'b1000000001101000: out_v[312] = 10'b0010101111;
    16'b0000010001101100: out_v[312] = 10'b0110011011;
    16'b0000000000001100: out_v[312] = 10'b1011010101;
    16'b0000010000100000: out_v[312] = 10'b1011101001;
    16'b0000000001001001: out_v[312] = 10'b1110101111;
    16'b0000010000101101: out_v[312] = 10'b0001011001;
    16'b1000000000101101: out_v[312] = 10'b1010100010;
    16'b0000000000001101: out_v[312] = 10'b0011001111;
    16'b0000010001001101: out_v[312] = 10'b1001110010;
    16'b0010000001000000: out_v[312] = 10'b0001000111;
    16'b0000000001001101: out_v[312] = 10'b1011011101;
    16'b0000010000001101: out_v[312] = 10'b1011010111;
    16'b1000010001100000: out_v[312] = 10'b0100010110;
    16'b1000000000100101: out_v[312] = 10'b1111100010;
    16'b0000000001000001: out_v[312] = 10'b1011110111;
    16'b0000010000100101: out_v[312] = 10'b0100011110;
    16'b0000010000101000: out_v[312] = 10'b0101100001;
    16'b0010010001000000: out_v[312] = 10'b0110111011;
    16'b1000010000101101: out_v[312] = 10'b0001101110;
    16'b0000000001001100: out_v[312] = 10'b1100100000;
    16'b0000000001100000: out_v[312] = 10'b0100011100;
    16'b0100010001100000: out_v[312] = 10'b0000011001;
    16'b0000000000100000: out_v[312] = 10'b0001010000;
    16'b1100010001101000: out_v[312] = 10'b1110011011;
    16'b1100000001000000: out_v[312] = 10'b1011001011;
    16'b0100010000100101: out_v[312] = 10'b1000010011;
    16'b0100010000100000: out_v[312] = 10'b0111001011;
    16'b0000010000100001: out_v[312] = 10'b0111110011;
    16'b0100010001101000: out_v[312] = 10'b1000011111;
    16'b0100010000101001: out_v[312] = 10'b1011011111;
    16'b1101000000100101: out_v[312] = 10'b1000111001;
    16'b0100000000101101: out_v[312] = 10'b1011011110;
    16'b0000000000100101: out_v[312] = 10'b0110001100;
    16'b1100000001100000: out_v[312] = 10'b1010001011;
    16'b0100010001100001: out_v[312] = 10'b1010000001;
    16'b0000010100101101: out_v[312] = 10'b1000011001;
    16'b1100000001001000: out_v[312] = 10'b0011111001;
    16'b0100000001100000: out_v[312] = 10'b1111001001;
    16'b0000010000101001: out_v[312] = 10'b1111010001;
    16'b0100010000100001: out_v[312] = 10'b1101110010;
    16'b0000010001100101: out_v[312] = 10'b0000111101;
    16'b0100000001101000: out_v[312] = 10'b0011001101;
    16'b1100010001100000: out_v[312] = 10'b0110010110;
    16'b0100010100101001: out_v[312] = 10'b1010110010;
    16'b0100000000001000: out_v[312] = 10'b1000101110;
    16'b0100010100100001: out_v[312] = 10'b1011110111;
    16'b0100000000000000: out_v[312] = 10'b0011011010;
    16'b1100000000101101: out_v[312] = 10'b1010111010;
    16'b1000010100101001: out_v[312] = 10'b1111100101;
    16'b0000000100101001: out_v[312] = 10'b1110110011;
    16'b0100000000001001: out_v[312] = 10'b0100010011;
    16'b0000000100000000: out_v[312] = 10'b0011010001;
    16'b0100000000100100: out_v[312] = 10'b1101010010;
    16'b0100000000001101: out_v[312] = 10'b1111110001;
    16'b1100010100101001: out_v[312] = 10'b0001110110;
    16'b0000000100100000: out_v[312] = 10'b0110110011;
    16'b0100000000001100: out_v[312] = 10'b1111001000;
    16'b0100000100101001: out_v[312] = 10'b0101100111;
    16'b0000010100101001: out_v[312] = 10'b1010000100;
    16'b1100000100101101: out_v[312] = 10'b0110110110;
    16'b0000010100100000: out_v[312] = 10'b1011100011;
    16'b0100000000101001: out_v[312] = 10'b1101110111;
    16'b0100000100101101: out_v[312] = 10'b0000111100;
    16'b1100000000101100: out_v[312] = 10'b0100111010;
    16'b0100000000100001: out_v[312] = 10'b1101010011;
    16'b0100000000000001: out_v[312] = 10'b1000111000;
    16'b0100010100101101: out_v[312] = 10'b1110000000;
    16'b0000010100101000: out_v[312] = 10'b1111011001;
    16'b1000010100101000: out_v[312] = 10'b0111010010;
    16'b1000000100101000: out_v[312] = 10'b0000111010;
    16'b0000000100101000: out_v[312] = 10'b0010110111;
    16'b1100000000101000: out_v[312] = 10'b0100111001;
    16'b0100010100101000: out_v[312] = 10'b0011001111;
    16'b1100000000100000: out_v[312] = 10'b1010011001;
    16'b1100000100101001: out_v[312] = 10'b0111110111;
    16'b0100000000000101: out_v[312] = 10'b1111000001;
    16'b1000000100101001: out_v[312] = 10'b1110011011;
    16'b0100000000100101: out_v[312] = 10'b0000100010;
    16'b1100000000100100: out_v[312] = 10'b0011011001;
    16'b0100010100100000: out_v[312] = 10'b0100111111;
    16'b1100000100100101: out_v[312] = 10'b0010010011;
    16'b0100100000001000: out_v[312] = 10'b1011100110;
    16'b0000100000001000: out_v[312] = 10'b1110110000;
    16'b1100000000000101: out_v[312] = 10'b1101100100;
    16'b0100010100100101: out_v[312] = 10'b1100100101;
    16'b0100100000001101: out_v[312] = 10'b1000100110;
    16'b1100000000100101: out_v[312] = 10'b0000111111;
    16'b0100100000001100: out_v[312] = 10'b0011001100;
    16'b0100010001100101: out_v[312] = 10'b0001010011;
    16'b0100100000101000: out_v[312] = 10'b1000100111;
    16'b0100110100101101: out_v[312] = 10'b0101110000;
    16'b1100010001100101: out_v[312] = 10'b1011000111;
    16'b1110000100000101: out_v[312] = 10'b1011100000;
    16'b1100000001000001: out_v[312] = 10'b1001100001;
    16'b0000010000100100: out_v[312] = 10'b0000101100;
    16'b0100010001100100: out_v[312] = 10'b1111101010;
    16'b1100010001100100: out_v[312] = 10'b1100111110;
    16'b1100010101100101: out_v[312] = 10'b1011011100;
    16'b1100000001100100: out_v[312] = 10'b1111001000;
    16'b1100000001000101: out_v[312] = 10'b1111010001;
    16'b1110010101100101: out_v[312] = 10'b0111011000;
    16'b1100000001000100: out_v[312] = 10'b1111001011;
    16'b1100010101000101: out_v[312] = 10'b0100110111;
    16'b1100010001000100: out_v[312] = 10'b1010110011;
    16'b1100010001000101: out_v[312] = 10'b1011111011;
    16'b0100000001100100: out_v[312] = 10'b0011101010;
    16'b1100000001100101: out_v[312] = 10'b1111110001;
    16'b1100010000000100: out_v[312] = 10'b1100000010;
    16'b1100010000000000: out_v[312] = 10'b0101010011;
    16'b1100010000000101: out_v[312] = 10'b0111110011;
    16'b0000010001100100: out_v[312] = 10'b1110111000;
    16'b1100000000000100: out_v[312] = 10'b1100101011;
    16'b1000000101000001: out_v[312] = 10'b1011111110;
    16'b0001010000100101: out_v[312] = 10'b1111100110;
    16'b0100000100001000: out_v[312] = 10'b0111100011;
    16'b0000000100101101: out_v[312] = 10'b0110100010;
    16'b0001000100101101: out_v[312] = 10'b0101011111;
    16'b0101010100101101: out_v[312] = 10'b0101011011;
    16'b0100000100001101: out_v[312] = 10'b0111110110;
    16'b0001000000101101: out_v[312] = 10'b0011100001;
    16'b1001010100101101: out_v[312] = 10'b1011111000;
    16'b0000000100001101: out_v[312] = 10'b1000000110;
    16'b0000010100100101: out_v[312] = 10'b1001001110;
    16'b0001010100101101: out_v[312] = 10'b1101001011;
    16'b0001010000101101: out_v[312] = 10'b1011010110;
    16'b0001000000001101: out_v[312] = 10'b1001110110;
    16'b0000000100100101: out_v[312] = 10'b1001110111;
    16'b0000000100000101: out_v[312] = 10'b0010001110;
    16'b1000000100101101: out_v[312] = 10'b0111101001;
    16'b0100000100101100: out_v[312] = 10'b0100101110;
    16'b0100000100101000: out_v[312] = 10'b0011000111;
    16'b0100010000001101: out_v[312] = 10'b1101011000;
    16'b0100100000000101: out_v[312] = 10'b1101001011;
    16'b0100010100001101: out_v[312] = 10'b0100110011;
    16'b0100010001101001: out_v[312] = 10'b0111101100;
    16'b0100000100100101: out_v[312] = 10'b1101001111;
    16'b0000010100100001: out_v[312] = 10'b1101001010;
    16'b0100000100000101: out_v[312] = 10'b1100001000;
    default: out_v[312] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000100000001000: out_v[313] = 10'b1101100001;
    16'b0100110100011000: out_v[313] = 10'b0100000101;
    16'b0100100100011000: out_v[313] = 10'b1111001001;
    16'b0100010110011000: out_v[313] = 10'b0011110111;
    16'b0100010010011000: out_v[313] = 10'b1001001011;
    16'b0100100100010000: out_v[313] = 10'b0011101011;
    16'b0000100000010000: out_v[313] = 10'b0001011010;
    16'b0000110000001000: out_v[313] = 10'b1001011000;
    16'b0100110010011000: out_v[313] = 10'b1100110011;
    16'b0100000100011000: out_v[313] = 10'b0111011011;
    16'b0000110000011000: out_v[313] = 10'b0001101111;
    16'b0000100000000000: out_v[313] = 10'b0010111100;
    16'b0100000100010000: out_v[313] = 10'b1111100110;
    16'b0000110010011000: out_v[313] = 10'b0010111001;
    16'b0100000110010000: out_v[313] = 10'b0111000111;
    16'b0100110000011000: out_v[313] = 10'b0010110111;
    16'b0100000110011000: out_v[313] = 10'b1001100111;
    16'b0000100000011000: out_v[313] = 10'b1000100110;
    16'b0100010110001000: out_v[313] = 10'b1001010111;
    16'b0000110010001000: out_v[313] = 10'b0110010011;
    16'b0100100100001000: out_v[313] = 10'b1001100010;
    16'b0100110110011000: out_v[313] = 10'b0001011011;
    16'b0000110100011000: out_v[313] = 10'b0010101010;
    16'b0100010100001000: out_v[313] = 10'b0110000011;
    16'b0000100010001000: out_v[313] = 10'b1101000001;
    16'b0100000010011000: out_v[313] = 10'b0010111101;
    16'b0100100000010000: out_v[313] = 10'b1000111011;
    16'b0100010100011000: out_v[313] = 10'b0010000101;
    16'b0000010010011000: out_v[313] = 10'b0100110011;
    16'b0100100110011000: out_v[313] = 10'b0001001010;
    16'b0000100100001000: out_v[313] = 10'b0111100010;
    16'b0100100100000000: out_v[313] = 10'b0100100001;
    16'b0000110100001000: out_v[313] = 10'b1011000011;
    16'b0100110100001000: out_v[313] = 10'b1011001000;
    16'b0100100000011000: out_v[313] = 10'b0010111110;
    16'b0000110000000000: out_v[313] = 10'b1101101100;
    16'b0000010110001000: out_v[313] = 10'b1010101010;
    16'b0000010010001000: out_v[313] = 10'b1011110000;
    16'b0000000000000000: out_v[313] = 10'b0010010110;
    16'b0000010010000000: out_v[313] = 10'b1001100111;
    16'b0000100010000000: out_v[313] = 10'b1101000010;
    16'b0000110010000000: out_v[313] = 10'b0110000111;
    16'b0000000010000000: out_v[313] = 10'b0011111100;
    16'b0000010100001000: out_v[313] = 10'b0100101011;
    16'b0000010110000000: out_v[313] = 10'b0011100000;
    16'b0100000110011001: out_v[313] = 10'b1011110010;
    16'b0000110110001000: out_v[313] = 10'b0101011110;
    16'b0000010110001001: out_v[313] = 10'b1010110100;
    16'b0100010110001001: out_v[313] = 10'b1101011100;
    16'b0000000110001000: out_v[313] = 10'b1001100101;
    16'b0000010000001001: out_v[313] = 10'b1010101101;
    16'b0100010010001000: out_v[313] = 10'b0000100110;
    16'b0100000100000000: out_v[313] = 10'b0110110011;
    16'b0100000110001000: out_v[313] = 10'b0011101110;
    16'b0100000010010000: out_v[313] = 10'b0111010011;
    16'b0100110110001000: out_v[313] = 10'b1001101000;
    16'b0100010010001001: out_v[313] = 10'b0110011001;
    16'b0100010010011001: out_v[313] = 10'b1100000111;
    16'b0100000010001000: out_v[313] = 10'b1000111010;
    16'b0100000110000001: out_v[313] = 10'b0111001110;
    16'b0100010000011000: out_v[313] = 10'b1111110110;
    16'b0000000110000000: out_v[313] = 10'b1110111000;
    16'b0100010000001000: out_v[313] = 10'b1001110100;
    16'b0100000110000000: out_v[313] = 10'b0000101100;
    16'b0000010000000000: out_v[313] = 10'b1101010000;
    16'b0100010010000000: out_v[313] = 10'b1000101110;
    16'b0000010010001001: out_v[313] = 10'b1110110101;
    16'b0100000110001001: out_v[313] = 10'b1101111100;
    16'b0000010010000001: out_v[313] = 10'b1101010110;
    16'b0100000110010001: out_v[313] = 10'b1010011010;
    16'b0000010000001000: out_v[313] = 10'b1110001001;
    16'b0100000010000000: out_v[313] = 10'b1110111000;
    16'b0100000100001000: out_v[313] = 10'b0100010101;
    16'b0100010110011001: out_v[313] = 10'b0100000011;
    16'b0000110100000000: out_v[313] = 10'b0111100000;
    16'b0000100100000000: out_v[313] = 10'b0010111000;
    16'b0100110100000000: out_v[313] = 10'b0011001100;
    16'b0000000100001000: out_v[313] = 10'b0111000010;
    16'b0000000100000000: out_v[313] = 10'b1100100001;
    16'b0100110000001000: out_v[313] = 10'b1010011011;
    16'b0000010000010000: out_v[313] = 10'b0111110000;
    16'b0000010000011000: out_v[313] = 10'b0011011000;
    16'b0000000010010000: out_v[313] = 10'b0101100000;
    16'b0000000010011000: out_v[313] = 10'b1100110000;
    16'b0000000000011000: out_v[313] = 10'b1110000101;
    16'b0000000110010000: out_v[313] = 10'b0001011111;
    16'b0000000000001000: out_v[313] = 10'b1100101011;
    16'b0000100010010000: out_v[313] = 10'b0100110010;
    16'b0000000000010000: out_v[313] = 10'b0000010110;
    16'b0100000000010000: out_v[313] = 10'b1111010110;
    16'b0000100100010000: out_v[313] = 10'b1100101010;
    16'b0100100000000000: out_v[313] = 10'b0000110011;
    16'b0000001000000000: out_v[313] = 10'b1011111000;
    16'b0000000010000001: out_v[313] = 10'b0011100000;
    16'b0000001010000001: out_v[313] = 10'b0011100011;
    16'b0000000010010001: out_v[313] = 10'b0110111011;
    16'b0000001010010001: out_v[313] = 10'b1111111101;
    16'b0000010010010000: out_v[313] = 10'b1101001101;
    16'b0000000000000001: out_v[313] = 10'b1101110000;
    16'b0100000010010001: out_v[313] = 10'b0001110110;
    16'b0100001010010001: out_v[313] = 10'b0101110010;
    16'b0100001010010000: out_v[313] = 10'b0011010010;
    16'b0000001010010000: out_v[313] = 10'b0111101011;
    16'b0000001010000000: out_v[313] = 10'b1111011101;
    16'b0100001010000000: out_v[313] = 10'b1111110011;
    16'b0000000000010001: out_v[313] = 10'b1011100100;
    16'b0000000010001000: out_v[313] = 10'b1010100001;
    16'b0000110000010000: out_v[313] = 10'b1010001101;
    16'b0000100110001000: out_v[313] = 10'b0001101111;
    16'b0000100110000000: out_v[313] = 10'b1100100110;
    16'b0000100010011000: out_v[313] = 10'b1000010010;
    default: out_v[313] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000100000000100: out_v[314] = 10'b0100011101;
    16'b1000000000000100: out_v[314] = 10'b1110100011;
    16'b1000000100010101: out_v[314] = 10'b1111001011;
    16'b1000000110000101: out_v[314] = 10'b1011101010;
    16'b0000000000000000: out_v[314] = 10'b0001100000;
    16'b1000000110010100: out_v[314] = 10'b0101001111;
    16'b1000000100000100: out_v[314] = 10'b0010011110;
    16'b1000000100000001: out_v[314] = 10'b0111011101;
    16'b1000000110000100: out_v[314] = 10'b0101001001;
    16'b1000000000000000: out_v[314] = 10'b1100011101;
    16'b0000100000010100: out_v[314] = 10'b1010100110;
    16'b1000000100000101: out_v[314] = 10'b0110011000;
    16'b0000000000010100: out_v[314] = 10'b0111011100;
    16'b0000000000000100: out_v[314] = 10'b1100100000;
    16'b0000000000000001: out_v[314] = 10'b0100100001;
    16'b1000000110000000: out_v[314] = 10'b0111001001;
    16'b1000000001000100: out_v[314] = 10'b1000101011;
    16'b1000000000010100: out_v[314] = 10'b0110011101;
    16'b1000000001000000: out_v[314] = 10'b1111011011;
    16'b1000000000000001: out_v[314] = 10'b1100011110;
    16'b0000000100000101: out_v[314] = 10'b1111100011;
    16'b1000000110000001: out_v[314] = 10'b0101111011;
    16'b0000000001000100: out_v[314] = 10'b0011110010;
    16'b1000000111000000: out_v[314] = 10'b0110011111;
    16'b1000000100010100: out_v[314] = 10'b1010000111;
    16'b0000000111000100: out_v[314] = 10'b0111111010;
    16'b1000100100010101: out_v[314] = 10'b1110010011;
    16'b1000000100000000: out_v[314] = 10'b1110010111;
    16'b0000000100010101: out_v[314] = 10'b1011000101;
    16'b1000000111000100: out_v[314] = 10'b1001001010;
    16'b0000000100000100: out_v[314] = 10'b1111100110;
    16'b1000100110010100: out_v[314] = 10'b0110110011;
    16'b1000000110010101: out_v[314] = 10'b0101001001;
    16'b0000000100000001: out_v[314] = 10'b1000100110;
    16'b0000000100000000: out_v[314] = 10'b1001110110;
    16'b0000100001010100: out_v[314] = 10'b1010001101;
    16'b0000100001000100: out_v[314] = 10'b0100011111;
    16'b0000100100010101: out_v[314] = 10'b0000001011;
    16'b0000000000010000: out_v[314] = 10'b0110011111;
    16'b0000100000010101: out_v[314] = 10'b0010001011;
    16'b0000000001010000: out_v[314] = 10'b1100001011;
    16'b0000010001010000: out_v[314] = 10'b1110101101;
    16'b0000000001010100: out_v[314] = 10'b0110001100;
    16'b0000100100000101: out_v[314] = 10'b1000010111;
    16'b0000110000000100: out_v[314] = 10'b1011000110;
    16'b0000100001000101: out_v[314] = 10'b1101011011;
    16'b0000000101000001: out_v[314] = 10'b0010100100;
    16'b0000100000000101: out_v[314] = 10'b0010011010;
    16'b0000000001000000: out_v[314] = 10'b0001101010;
    16'b0000110001010100: out_v[314] = 10'b0111011111;
    16'b0000100001010101: out_v[314] = 10'b1001101100;
    16'b0000100100010100: out_v[314] = 10'b1010001010;
    16'b0000100100000100: out_v[314] = 10'b0000011001;
    16'b0000100101010100: out_v[314] = 10'b0001011100;
    16'b0000110001000100: out_v[314] = 10'b0000010111;
    16'b0000010001010100: out_v[314] = 10'b0100110011;
    16'b0000010000010000: out_v[314] = 10'b0010101111;
    16'b0000000000000101: out_v[314] = 10'b1101110010;
    16'b0000110000010100: out_v[314] = 10'b1011111011;
    16'b0000100101000101: out_v[314] = 10'b1100000011;
    16'b0000100101000100: out_v[314] = 10'b0110001110;
    16'b0000100100000001: out_v[314] = 10'b1001111011;
    16'b0000000000010101: out_v[314] = 10'b1000111100;
    16'b0000100000000001: out_v[314] = 10'b0111011001;
    16'b0000100001010000: out_v[314] = 10'b1001110101;
    16'b0000100000000000: out_v[314] = 10'b1100011010;
    16'b0000100000010000: out_v[314] = 10'b1011100110;
    16'b0000000001010101: out_v[314] = 10'b0011001011;
    16'b0000100010000100: out_v[314] = 10'b0111010101;
    16'b0000100100000000: out_v[314] = 10'b0101111100;
    16'b0000000100010100: out_v[314] = 10'b1000101000;
    16'b0000000010000000: out_v[314] = 10'b1101011110;
    16'b0000100010010100: out_v[314] = 10'b1100010110;
    16'b0000100110000100: out_v[314] = 10'b0000111011;
    16'b0000000110000000: out_v[314] = 10'b1001010110;
    16'b1000100000010100: out_v[314] = 10'b1011110110;
    16'b0000000001000001: out_v[314] = 10'b1111100010;
    16'b0000000011000000: out_v[314] = 10'b0010100010;
    16'b0000010001000000: out_v[314] = 10'b1111000100;
    16'b0000010000000000: out_v[314] = 10'b1110001100;
    16'b1000100000000000: out_v[314] = 10'b1011000100;
    16'b0000110000000000: out_v[314] = 10'b1111101011;
    16'b0000101000000100: out_v[314] = 10'b1000001110;
    16'b0000101000010100: out_v[314] = 10'b0110101001;
    16'b0000001000000100: out_v[314] = 10'b1001000111;
    16'b0000001000010100: out_v[314] = 10'b0110100100;
    16'b0100100010010100: out_v[314] = 10'b0011110111;
    16'b0000101010010100: out_v[314] = 10'b1101100011;
    16'b1000100000000100: out_v[314] = 10'b1001000110;
    16'b0000100011010100: out_v[314] = 10'b1110010111;
    default: out_v[314] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000001000000000: out_v[315] = 10'b1010111110;
    16'b0101001000001000: out_v[315] = 10'b0111000011;
    16'b0000001010001000: out_v[315] = 10'b1100011011;
    16'b0001001100001000: out_v[315] = 10'b1100000001;
    16'b0001001010001000: out_v[315] = 10'b0001011110;
    16'b0001001000001000: out_v[315] = 10'b0101011101;
    16'b0000001000001000: out_v[315] = 10'b1000100111;
    16'b0101001000000000: out_v[315] = 10'b0101101011;
    16'b0101000010001000: out_v[315] = 10'b1100011011;
    16'b0001001010001010: out_v[315] = 10'b1000110010;
    16'b0100001000000000: out_v[315] = 10'b1010101010;
    16'b0100001000001000: out_v[315] = 10'b1001110100;
    16'b0101001100001000: out_v[315] = 10'b1011100001;
    16'b0001101100001000: out_v[315] = 10'b0100011011;
    16'b0101001110001000: out_v[315] = 10'b1011000111;
    16'b0101001010001000: out_v[315] = 10'b0100101101;
    16'b0101101000001000: out_v[315] = 10'b0011101111;
    16'b0101001010001010: out_v[315] = 10'b0001000011;
    16'b0101000000001000: out_v[315] = 10'b0110101011;
    16'b0001000010001010: out_v[315] = 10'b0110000101;
    16'b0001001000000000: out_v[315] = 10'b1011000101;
    16'b0000001010001010: out_v[315] = 10'b0000101101;
    16'b1000001000000000: out_v[315] = 10'b0001010111;
    16'b0100101000001000: out_v[315] = 10'b0011111000;
    16'b1000000010001010: out_v[315] = 10'b1010111111;
    16'b1000001010000010: out_v[315] = 10'b1110011100;
    16'b0000001010000010: out_v[315] = 10'b0111100110;
    16'b1000000010000010: out_v[315] = 10'b1100011101;
    16'b1000000000000000: out_v[315] = 10'b1010010010;
    16'b1000001010000000: out_v[315] = 10'b0101111011;
    16'b0000000010000010: out_v[315] = 10'b0111000010;
    16'b1000000000000010: out_v[315] = 10'b1101000100;
    16'b1000000000001010: out_v[315] = 10'b0011011010;
    16'b1000000000001000: out_v[315] = 10'b1000111010;
    16'b1000001010001010: out_v[315] = 10'b0111000000;
    16'b1000000010000000: out_v[315] = 10'b0101011100;
    16'b0000100010000010: out_v[315] = 10'b1111100011;
    16'b0000001010000000: out_v[315] = 10'b0011001110;
    16'b1000001010001110: out_v[315] = 10'b1110101001;
    16'b1000000010001110: out_v[315] = 10'b0110011101;
    16'b1001000010001010: out_v[315] = 10'b0001000100;
    16'b1000001000000010: out_v[315] = 10'b1100001001;
    16'b1001001010001110: out_v[315] = 10'b1001110111;
    16'b1101000010001010: out_v[315] = 10'b1001100101;
    16'b1001000010001110: out_v[315] = 10'b0010100110;
    16'b0000000010001010: out_v[315] = 10'b1011100111;
    16'b1001001010001010: out_v[315] = 10'b1010110000;
    16'b1001000010000010: out_v[315] = 10'b0000010110;
    16'b1000001000001000: out_v[315] = 10'b0001000100;
    16'b1001000110001010: out_v[315] = 10'b0000000100;
    16'b1000001010001000: out_v[315] = 10'b0101111101;
    16'b1001000010001000: out_v[315] = 10'b0011100110;
    16'b1000001000001010: out_v[315] = 10'b0101110100;
    16'b0001000010001110: out_v[315] = 10'b1011011111;
    16'b1101000110001010: out_v[315] = 10'b1101101110;
    16'b0000001010001110: out_v[315] = 10'b1011110011;
    16'b1000000010001000: out_v[315] = 10'b1101110001;
    16'b1000001000001100: out_v[315] = 10'b0100100110;
    16'b1001000000001010: out_v[315] = 10'b0001010111;
    16'b0000000010001110: out_v[315] = 10'b1001100010;
    16'b1000001000001110: out_v[315] = 10'b1011000101;
    16'b1001000000000010: out_v[315] = 10'b0110000111;
    16'b0000001000000010: out_v[315] = 10'b0000111000;
    16'b0000101000000000: out_v[315] = 10'b1011100111;
    16'b0000101000001010: out_v[315] = 10'b0110011111;
    16'b0000101000001000: out_v[315] = 10'b0001001011;
    16'b0000101000000010: out_v[315] = 10'b1011111000;
    16'b0000100000000010: out_v[315] = 10'b0001111011;
    16'b0000000000000010: out_v[315] = 10'b0001011000;
    16'b0000100000000000: out_v[315] = 10'b0111001100;
    16'b0000001000001010: out_v[315] = 10'b0010101101;
    16'b0001001000001010: out_v[315] = 10'b0000101010;
    16'b0100101000000000: out_v[315] = 10'b1001110011;
    16'b0001001000001100: out_v[315] = 10'b0110011101;
    16'b0000000000000000: out_v[315] = 10'b1000011101;
    16'b0000001000001100: out_v[315] = 10'b1010100101;
    16'b1000100010000010: out_v[315] = 10'b1001101001;
    16'b1001001010000010: out_v[315] = 10'b0110010010;
    16'b1100001010000010: out_v[315] = 10'b0011111000;
    16'b1000100000000010: out_v[315] = 10'b0111010011;
    16'b1101001010000010: out_v[315] = 10'b0110111000;
    16'b1100000000000010: out_v[315] = 10'b1111101001;
    16'b1101000010000010: out_v[315] = 10'b0010010111;
    16'b1100000010000010: out_v[315] = 10'b0110101011;
    16'b0001001010000010: out_v[315] = 10'b0110010010;
    16'b0100001010000010: out_v[315] = 10'b1111000001;
    16'b0100000000000010: out_v[315] = 10'b0011011010;
    16'b1101000000000010: out_v[315] = 10'b1100111110;
    16'b1001100010000010: out_v[315] = 10'b0011001001;
    16'b0001000010001000: out_v[315] = 10'b0100011010;
    16'b1000101010000010: out_v[315] = 10'b0100110110;
    16'b1100001010001010: out_v[315] = 10'b1110110111;
    16'b1000000010000100: out_v[315] = 10'b1011000101;
    16'b1100000010000110: out_v[315] = 10'b1010101101;
    16'b1000000000000100: out_v[315] = 10'b0111011100;
    16'b0100000010000110: out_v[315] = 10'b0110100011;
    16'b1000001010000110: out_v[315] = 10'b1001001011;
    16'b0100000010001010: out_v[315] = 10'b1111011010;
    16'b1101001010001010: out_v[315] = 10'b1011001101;
    16'b1100001010000110: out_v[315] = 10'b1011001100;
    16'b1100000010000000: out_v[315] = 10'b1111000011;
    16'b1100000010001010: out_v[315] = 10'b0100111011;
    16'b1100000010001110: out_v[315] = 10'b0110111111;
    16'b0000000010000110: out_v[315] = 10'b1101101110;
    16'b1000000010000110: out_v[315] = 10'b1111111101;
    16'b0100000010000010: out_v[315] = 10'b0011101011;
    16'b0101000010001010: out_v[315] = 10'b0101010110;
    16'b1100000010000100: out_v[315] = 10'b1111111011;
    16'b0000001011000010: out_v[315] = 10'b1001000111;
    16'b0000000011000010: out_v[315] = 10'b1101001001;
    16'b0000101010000010: out_v[315] = 10'b0100000101;
    16'b0000001011000000: out_v[315] = 10'b1110010111;
    16'b0000001001000000: out_v[315] = 10'b1101111100;
    16'b1000001011000010: out_v[315] = 10'b1000111010;
    16'b1000000011000010: out_v[315] = 10'b0111110001;
    16'b0100100000000000: out_v[315] = 10'b0010110010;
    16'b1001001000001010: out_v[315] = 10'b1101101001;
    16'b1000101000000000: out_v[315] = 10'b0111000111;
    16'b1000101000000010: out_v[315] = 10'b0101010110;
    16'b1000101010001010: out_v[315] = 10'b0101010100;
    16'b1000101000001010: out_v[315] = 10'b1011110111;
    16'b1000100000000000: out_v[315] = 10'b1101100100;
    default: out_v[315] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000001100000010: out_v[316] = 10'b1111010001;
    16'b0000001101000001: out_v[316] = 10'b0010110011;
    16'b1000001001100111: out_v[316] = 10'b1011100011;
    16'b1000001001100011: out_v[316] = 10'b0000110001;
    16'b0000001100000011: out_v[316] = 10'b1100011011;
    16'b0000001100000000: out_v[316] = 10'b0010110011;
    16'b1000001001100001: out_v[316] = 10'b0000000011;
    16'b1000000001100011: out_v[316] = 10'b1011011000;
    16'b0000000100000010: out_v[316] = 10'b0011011101;
    16'b0000001101100001: out_v[316] = 10'b1111111001;
    16'b1000000001100001: out_v[316] = 10'b0011000011;
    16'b1000001101100001: out_v[316] = 10'b1110100111;
    16'b0000000101000001: out_v[316] = 10'b1010000111;
    16'b0000001101000011: out_v[316] = 10'b1011001011;
    16'b0000001001000011: out_v[316] = 10'b1101100110;
    16'b0000000001000011: out_v[316] = 10'b1010011101;
    16'b1010001001100011: out_v[316] = 10'b0011100010;
    16'b1000001101100011: out_v[316] = 10'b0011010101;
    16'b1000001001000011: out_v[316] = 10'b0101111110;
    16'b0000001100000001: out_v[316] = 10'b0101100011;
    16'b0000000101100001: out_v[316] = 10'b1011011101;
    16'b0000001101000000: out_v[316] = 10'b0010111100;
    16'b0000000100000000: out_v[316] = 10'b1001100111;
    16'b0000001000000010: out_v[316] = 10'b1000000111;
    16'b1000000101100001: out_v[316] = 10'b0000000111;
    16'b1000001000100011: out_v[316] = 10'b1010011011;
    16'b0010001001000011: out_v[316] = 10'b1111010100;
    16'b0000001000000011: out_v[316] = 10'b1100001110;
    16'b1010001001100111: out_v[316] = 10'b1110101111;
    16'b1000001001100010: out_v[316] = 10'b0111011011;
    16'b0000001101100011: out_v[316] = 10'b1111100011;
    16'b0000000000010000: out_v[316] = 10'b1110001010;
    16'b0000000000010010: out_v[316] = 10'b1110000001;
    16'b0000000000000000: out_v[316] = 10'b1101011111;
    16'b0000000010010000: out_v[316] = 10'b0010001011;
    16'b0000000000000010: out_v[316] = 10'b1011110000;
    16'b0000001000010000: out_v[316] = 10'b0110001010;
    16'b0000000010010010: out_v[316] = 10'b1001001010;
    16'b0000000100010000: out_v[316] = 10'b0001000000;
    16'b0010000000010010: out_v[316] = 10'b1110100011;
    16'b0010000000010000: out_v[316] = 10'b1111100101;
    16'b0010000000000010: out_v[316] = 10'b0010110010;
    16'b0000000000010110: out_v[316] = 10'b1001101100;
    16'b0010000000000000: out_v[316] = 10'b0010010101;
    16'b0010000000010100: out_v[316] = 10'b1111000101;
    16'b0000000100010010: out_v[316] = 10'b1010111000;
    16'b1000001100110000: out_v[316] = 10'b1110000111;
    16'b0011000000010110: out_v[316] = 10'b1111111001;
    16'b0010000000010110: out_v[316] = 10'b0101100101;
    16'b0010000000000100: out_v[316] = 10'b0001111101;
    16'b0001000000010010: out_v[316] = 10'b0010111101;
    16'b0010000000000110: out_v[316] = 10'b1110010101;
    16'b0000001000000110: out_v[316] = 10'b1010100100;
    16'b0010001000010010: out_v[316] = 10'b0110110011;
    16'b0010001000010000: out_v[316] = 10'b1010010111;
    16'b0000001000110010: out_v[316] = 10'b0011001111;
    16'b0010001000000110: out_v[316] = 10'b1100110101;
    16'b0011000000010010: out_v[316] = 10'b1110111001;
    16'b0000001000010010: out_v[316] = 10'b0100001001;
    16'b1000001100110010: out_v[316] = 10'b0100110110;
    16'b0000001100010010: out_v[316] = 10'b1000010110;
    16'b0010001000010110: out_v[316] = 10'b1101100110;
    16'b0010001000000000: out_v[316] = 10'b1110110001;
    16'b0000001000000000: out_v[316] = 10'b1010010101;
    16'b0010001000000010: out_v[316] = 10'b1011101000;
    16'b0000001000110000: out_v[316] = 10'b0111111001;
    16'b0000000000010011: out_v[316] = 10'b0011010111;
    16'b0010000100010000: out_v[316] = 10'b0000001011;
    16'b0000001000100010: out_v[316] = 10'b1111000001;
    16'b0010000100010010: out_v[316] = 10'b0010101111;
    16'b0000000000000110: out_v[316] = 10'b1000010011;
    16'b0000000000010001: out_v[316] = 10'b0110000111;
    16'b1000001000110010: out_v[316] = 10'b0010001001;
    16'b1000001100111000: out_v[316] = 10'b1111100101;
    16'b0010000100000000: out_v[316] = 10'b1000000110;
    16'b0010000100010111: out_v[316] = 10'b0100011011;
    16'b0000001100010000: out_v[316] = 10'b1101011101;
    16'b0010000100000111: out_v[316] = 10'b0100110111;
    16'b0010001100010010: out_v[316] = 10'b0111111001;
    16'b0010000110010110: out_v[316] = 10'b0111000011;
    16'b0010000110010111: out_v[316] = 10'b1011110111;
    16'b0000000110010110: out_v[316] = 10'b1001101101;
    16'b0010000100000010: out_v[316] = 10'b0100011000;
    16'b0000000110010010: out_v[316] = 10'b1001111101;
    16'b0010000000000111: out_v[316] = 10'b1001111010;
    16'b0010000000000011: out_v[316] = 10'b0010101011;
    16'b0010000100010011: out_v[316] = 10'b1000100110;
    16'b0010000100010110: out_v[316] = 10'b0010101111;
    16'b0010000000000001: out_v[316] = 10'b0100111001;
    16'b0010000100000001: out_v[316] = 10'b1101100110;
    16'b0000000000000111: out_v[316] = 10'b1110100000;
    16'b0010000110000111: out_v[316] = 10'b1011011000;
    16'b0000000010010110: out_v[316] = 10'b0011011011;
    16'b0000000100010111: out_v[316] = 10'b0111001011;
    16'b0010000100000011: out_v[316] = 10'b0011000101;
    16'b0000000100000011: out_v[316] = 10'b1101001110;
    16'b0000000110010000: out_v[316] = 10'b0011010001;
    16'b0000000100010011: out_v[316] = 10'b1100110011;
    16'b0000001101010010: out_v[316] = 10'b0100110000;
    16'b0000001100010011: out_v[316] = 10'b0111010111;
    16'b0000001110010010: out_v[316] = 10'b0101001010;
    16'b1000001100010010: out_v[316] = 10'b0011111011;
    16'b0000000110000010: out_v[316] = 10'b1001100101;
    16'b0000001101010000: out_v[316] = 10'b1100111010;
    16'b0000000100010100: out_v[316] = 10'b0010111011;
    16'b0000000110000000: out_v[316] = 10'b1100100010;
    16'b1000001100010000: out_v[316] = 10'b0100011010;
    16'b1000001100010011: out_v[316] = 10'b0110011110;
    16'b0000000100010001: out_v[316] = 10'b1100111101;
    16'b0000001100010001: out_v[316] = 10'b0000110011;
    16'b0000000110010100: out_v[316] = 10'b0001110101;
    16'b1000000100010001: out_v[316] = 10'b1111111000;
    16'b1000001100010001: out_v[316] = 10'b0110111011;
    16'b0010000110010010: out_v[316] = 10'b1011011001;
    16'b0000000000100000: out_v[316] = 10'b1101110010;
    16'b0000000000000011: out_v[316] = 10'b1110100001;
    16'b1000000000100000: out_v[316] = 10'b0100110101;
    16'b0000000100110000: out_v[316] = 10'b0010111011;
    16'b0000001100110000: out_v[316] = 10'b1111110010;
    16'b0000000100100000: out_v[316] = 10'b1010010000;
    16'b0000000010000010: out_v[316] = 10'b1100000100;
    16'b0000000100000001: out_v[316] = 10'b1111100110;
    16'b0000010100010001: out_v[316] = 10'b1010101001;
    16'b0000010000010011: out_v[316] = 10'b1110111011;
    16'b0000010100000001: out_v[316] = 10'b0001000010;
    16'b0000010100010000: out_v[316] = 10'b1111001101;
    16'b0000010100000000: out_v[316] = 10'b1111010100;
    16'b0000010100010011: out_v[316] = 10'b1110010101;
    16'b0000001001010011: out_v[316] = 10'b1011100011;
    16'b0000010100000011: out_v[316] = 10'b1101011111;
    16'b0000001101010011: out_v[316] = 10'b1001000001;
    16'b0000001001000100: out_v[316] = 10'b1011000111;
    16'b0000000010000110: out_v[316] = 10'b0111110000;
    16'b0000001001000000: out_v[316] = 10'b0110110100;
    16'b0000000010000100: out_v[316] = 10'b0110100111;
    16'b0000000000000100: out_v[316] = 10'b0001011010;
    16'b0000001010000100: out_v[316] = 10'b0010001111;
    16'b0000001001000010: out_v[316] = 10'b0110011111;
    16'b0000001010000110: out_v[316] = 10'b1001110111;
    16'b0000000010000000: out_v[316] = 10'b0100110101;
    16'b0000001001000111: out_v[316] = 10'b0010110000;
    16'b0000001001000110: out_v[316] = 10'b1010110001;
    16'b0000001000000100: out_v[316] = 10'b0000100111;
    16'b0000001010000000: out_v[316] = 10'b1011100000;
    16'b0000001001000101: out_v[316] = 10'b1111101011;
    16'b0000000000010111: out_v[316] = 10'b1000011111;
    16'b0000001001010010: out_v[316] = 10'b0011011011;
    16'b0000001001010000: out_v[316] = 10'b0011100000;
    16'b0000001110010110: out_v[316] = 10'b0101111011;
    16'b0000000001010010: out_v[316] = 10'b0110011011;
    16'b0000001010010010: out_v[316] = 10'b0011011111;
    16'b0000001111010010: out_v[316] = 10'b0111110010;
    16'b0000001010000010: out_v[316] = 10'b1001100101;
    16'b0000001110000010: out_v[316] = 10'b0001111101;
    default: out_v[316] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1010000001000000: out_v[317] = 10'b1110001101;
    16'b1010000000000100: out_v[317] = 10'b0110110000;
    16'b1011010001000100: out_v[317] = 10'b1000101111;
    16'b1011000001000000: out_v[317] = 10'b0101011010;
    16'b1011000000000000: out_v[317] = 10'b0001010001;
    16'b0010000000000100: out_v[317] = 10'b0111001101;
    16'b1001000001000100: out_v[317] = 10'b0011101011;
    16'b1010010001000100: out_v[317] = 10'b0110000111;
    16'b1001000001000000: out_v[317] = 10'b0110001111;
    16'b1010000001000100: out_v[317] = 10'b1000001011;
    16'b1000000001000100: out_v[317] = 10'b1011011011;
    16'b1010010001000000: out_v[317] = 10'b1011111000;
    16'b1011000001000100: out_v[317] = 10'b0101110100;
    16'b1000000001000000: out_v[317] = 10'b1011001000;
    16'b0010010001000100: out_v[317] = 10'b0011011010;
    16'b0010000000000000: out_v[317] = 10'b0011100100;
    16'b1011010001000000: out_v[317] = 10'b0011110000;
    16'b1001010001000100: out_v[317] = 10'b1010101110;
    16'b1000000000000100: out_v[317] = 10'b0101010010;
    16'b1010000000000000: out_v[317] = 10'b1100010011;
    16'b0010000001000100: out_v[317] = 10'b0100010011;
    16'b1000010001000100: out_v[317] = 10'b1110100010;
    16'b0000000000000100: out_v[317] = 10'b0011001101;
    16'b1001000000000000: out_v[317] = 10'b0100011011;
    16'b1000000000000000: out_v[317] = 10'b0000110100;
    16'b1110010001000100: out_v[317] = 10'b0010101101;
    16'b1010010000000000: out_v[317] = 10'b1100000101;
    16'b0000000001000000: out_v[317] = 10'b0100110000;
    16'b0000000000000000: out_v[317] = 10'b1010100010;
    16'b0000010001000000: out_v[317] = 10'b1101100111;
    16'b0000010000000000: out_v[317] = 10'b0100110100;
    16'b1000010001000000: out_v[317] = 10'b0101100101;
    16'b0010000000011000: out_v[317] = 10'b1001010010;
    16'b0010000000001000: out_v[317] = 10'b0111010011;
    16'b0010010001000000: out_v[317] = 10'b0000011101;
    16'b0110010001000000: out_v[317] = 10'b0010111011;
    16'b1111010001000100: out_v[317] = 10'b0111110011;
    16'b1111010001000000: out_v[317] = 10'b1000011100;
    16'b1110010001000000: out_v[317] = 10'b0010110101;
    16'b1101010000000000: out_v[317] = 10'b1011010110;
    16'b1011010000000000: out_v[317] = 10'b1110001111;
    16'b1111010000000000: out_v[317] = 10'b0000011100;
    16'b1001010000000000: out_v[317] = 10'b1111010110;
    16'b0111010000000000: out_v[317] = 10'b0110111110;
    16'b1010010001000010: out_v[317] = 10'b0010001111;
    16'b1110010000000000: out_v[317] = 10'b0010001100;
    16'b1001010001000000: out_v[317] = 10'b1111100110;
    16'b0011010000000000: out_v[317] = 10'b1110101100;
    16'b1011000001000001: out_v[317] = 10'b0000000110;
    16'b1011010001000010: out_v[317] = 10'b0000011101;
    16'b1100010001000000: out_v[317] = 10'b1110101001;
    16'b0010000001000000: out_v[317] = 10'b0101110010;
    16'b1011000001011000: out_v[317] = 10'b0001000111;
    16'b0110010001000100: out_v[317] = 10'b0011011010;
    16'b1011010001000001: out_v[317] = 10'b1111000100;
    16'b1111010000000100: out_v[317] = 10'b0011011111;
    16'b1001000001000001: out_v[317] = 10'b1011101000;
    16'b1000000001000001: out_v[317] = 10'b0111011011;
    16'b0000000001000100: out_v[317] = 10'b0100011110;
    16'b1001010001000001: out_v[317] = 10'b1010011001;
    16'b0000010001000100: out_v[317] = 10'b1101011010;
    16'b1000010000000000: out_v[317] = 10'b0111001101;
    16'b0000000000010000: out_v[317] = 10'b0101010001;
    16'b0000000000011000: out_v[317] = 10'b1001100100;
    16'b0000000000001000: out_v[317] = 10'b1011110110;
    16'b0001000000000000: out_v[317] = 10'b1111001110;
    16'b1010000001011000: out_v[317] = 10'b1110110100;
    16'b1010000000011000: out_v[317] = 10'b0101101000;
    16'b1000000001011000: out_v[317] = 10'b0110110000;
    16'b1010000000010000: out_v[317] = 10'b1100001101;
    16'b1000000000010000: out_v[317] = 10'b1001101110;
    16'b1001000001001000: out_v[317] = 10'b1000110010;
    16'b1000000000011000: out_v[317] = 10'b0111101110;
    16'b1010000001010000: out_v[317] = 10'b1110110000;
    16'b0010000000010000: out_v[317] = 10'b1010100011;
    16'b1000000001001000: out_v[317] = 10'b0111011011;
    16'b1000000001010000: out_v[317] = 10'b0010110110;
    16'b1001000001011000: out_v[317] = 10'b0100110110;
    16'b0000001000000000: out_v[317] = 10'b1010101111;
    16'b0011000001000000: out_v[317] = 10'b0100100000;
    16'b0110010000000100: out_v[317] = 10'b0001000010;
    16'b0001000001000000: out_v[317] = 10'b1111100110;
    16'b0010010000000100: out_v[317] = 10'b1001011110;
    16'b0100010000000000: out_v[317] = 10'b1101100010;
    16'b0010010000000000: out_v[317] = 10'b1101110111;
    16'b0011010001000100: out_v[317] = 10'b1111000110;
    16'b0100010000000100: out_v[317] = 10'b0011111011;
    16'b0100010001000000: out_v[317] = 10'b0110010111;
    16'b0011000001000100: out_v[317] = 10'b1101010011;
    16'b0110010000000000: out_v[317] = 10'b1111000010;
    16'b0110000000000100: out_v[317] = 10'b0111011110;
    16'b0000100000100000: out_v[317] = 10'b1110111101;
    default: out_v[317] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010000000000111: out_v[318] = 10'b0101011011;
    16'b0010000000000110: out_v[318] = 10'b0111011011;
    16'b0000001000010111: out_v[318] = 10'b0010110110;
    16'b0001000000011101: out_v[318] = 10'b0110111110;
    16'b0000000000010001: out_v[318] = 10'b1001101011;
    16'b0100000000000100: out_v[318] = 10'b1110100101;
    16'b0010001000010111: out_v[318] = 10'b0100011011;
    16'b0100000000000110: out_v[318] = 10'b1000100111;
    16'b0000000000010101: out_v[318] = 10'b0101110101;
    16'b0000000000000100: out_v[318] = 10'b0010100011;
    16'b0100000000010101: out_v[318] = 10'b0100010101;
    16'b0110000000000100: out_v[318] = 10'b1011100100;
    16'b0010000000000000: out_v[318] = 10'b0110010110;
    16'b0010000000010111: out_v[318] = 10'b0010110010;
    16'b0010000000010101: out_v[318] = 10'b0101110100;
    16'b0110000000000000: out_v[318] = 10'b1001001011;
    16'b0010000000010001: out_v[318] = 10'b1110100100;
    16'b0010000000000101: out_v[318] = 10'b1101001111;
    16'b0010000000000100: out_v[318] = 10'b1010110010;
    16'b0000000000000110: out_v[318] = 10'b1100011101;
    16'b0000000000000101: out_v[318] = 10'b1100000111;
    16'b0011100000011101: out_v[318] = 10'b0001011111;
    16'b0000000000010111: out_v[318] = 10'b1001100000;
    16'b0100000000010111: out_v[318] = 10'b1110101101;
    16'b0000000000000111: out_v[318] = 10'b1010100101;
    16'b0001000000010101: out_v[318] = 10'b1111101000;
    16'b0011100100011101: out_v[318] = 10'b1111010111;
    16'b0100000000000000: out_v[318] = 10'b1100010111;
    16'b0000001000010101: out_v[318] = 10'b0000011010;
    16'b0010001000010101: out_v[318] = 10'b1011010100;
    16'b0100000000010110: out_v[318] = 10'b1010111111;
    16'b0110000000010001: out_v[318] = 10'b0100111001;
    16'b0000000000000000: out_v[318] = 10'b0001011111;
    16'b0100000000000101: out_v[318] = 10'b1011000010;
    16'b0010000000010011: out_v[318] = 10'b1110100101;
    16'b0110000000010101: out_v[318] = 10'b1111011110;
    16'b0110000000010111: out_v[318] = 10'b1110110011;
    16'b0011100000010101: out_v[318] = 10'b1100110101;
    16'b0100001000010111: out_v[318] = 10'b1001011011;
    16'b0100001000010101: out_v[318] = 10'b0011000111;
    16'b0100000000010001: out_v[318] = 10'b0100110011;
    16'b0000000000010000: out_v[318] = 10'b0110001011;
    16'b0000000000010100: out_v[318] = 10'b1011010010;
    16'b0010000000010000: out_v[318] = 10'b0011001010;
    16'b0000001000010001: out_v[318] = 10'b0010110100;
    16'b0000001000010000: out_v[318] = 10'b1110000010;
    16'b0100001000010001: out_v[318] = 10'b1100010000;
    16'b0010001000010000: out_v[318] = 10'b0101001011;
    16'b0000001000010100: out_v[318] = 10'b1001011100;
    16'b0110001000010101: out_v[318] = 10'b0101000111;
    16'b0000001000010011: out_v[318] = 10'b0000010110;
    16'b0001101100010101: out_v[318] = 10'b0111010111;
    16'b0000101000010101: out_v[318] = 10'b1011000011;
    16'b0000001000000101: out_v[318] = 10'b0111011000;
    16'b0001001000010001: out_v[318] = 10'b1100010110;
    16'b0001101100010011: out_v[318] = 10'b0111111011;
    16'b0001001000010101: out_v[318] = 10'b1001001101;
    16'b0000000000000010: out_v[318] = 10'b0111000110;
    16'b0000001000000000: out_v[318] = 10'b1001101001;
    16'b0001101100010111: out_v[318] = 10'b1000101110;
    16'b0001101000010101: out_v[318] = 10'b1011011000;
    16'b0001001000010011: out_v[318] = 10'b1110111011;
    16'b0000001000000111: out_v[318] = 10'b1111101001;
    16'b0000101000010001: out_v[318] = 10'b1100110010;
    16'b0100101000010101: out_v[318] = 10'b1110111001;
    16'b0000001000000011: out_v[318] = 10'b0011010000;
    16'b0001001100010101: out_v[318] = 10'b1101101101;
    16'b0000101000010111: out_v[318] = 10'b1011010010;
    16'b0100001000000101: out_v[318] = 10'b1001000101;
    16'b0001001100010111: out_v[318] = 10'b1110100111;
    16'b0000001000000001: out_v[318] = 10'b1000011100;
    16'b0010101000010101: out_v[318] = 10'b1111110011;
    16'b0000101100010101: out_v[318] = 10'b1111111111;
    16'b0010001000010001: out_v[318] = 10'b0101010111;
    16'b0001101100010001: out_v[318] = 10'b1001100110;
    16'b0000000000010011: out_v[318] = 10'b1000101011;
    16'b0000101000010011: out_v[318] = 10'b0010101111;
    16'b0000001000000010: out_v[318] = 10'b0001100100;
    16'b0000001000000100: out_v[318] = 10'b0110100000;
    16'b0110001000010001: out_v[318] = 10'b0101001011;
    16'b0110000000010000: out_v[318] = 10'b1111110111;
    16'b0110001000010011: out_v[318] = 10'b1010001010;
    16'b0010000000010010: out_v[318] = 10'b1101011000;
    16'b0100001000010011: out_v[318] = 10'b0111010010;
    16'b0010001000010011: out_v[318] = 10'b0011010111;
    16'b0010001000010100: out_v[318] = 10'b1111011001;
    16'b0100001000000001: out_v[318] = 10'b0101000011;
    16'b0010001000000000: out_v[318] = 10'b1110100010;
    16'b0010000000010100: out_v[318] = 10'b1101001000;
    16'b0110001000000101: out_v[318] = 10'b1101110111;
    16'b0110001000000001: out_v[318] = 10'b0000001011;
    16'b0110001000010111: out_v[318] = 10'b1011111000;
    16'b0010001000000100: out_v[318] = 10'b0000100111;
    16'b0110001000000000: out_v[318] = 10'b1000110110;
    16'b0110000000010011: out_v[318] = 10'b0011100010;
    16'b0110001000000011: out_v[318] = 10'b0011011011;
    16'b0000001000010010: out_v[318] = 10'b1011100001;
    16'b0010001000000011: out_v[318] = 10'b1110011110;
    16'b0000001000011011: out_v[318] = 10'b1000100011;
    16'b0010001000000010: out_v[318] = 10'b1000101100;
    16'b0000001000000110: out_v[318] = 10'b0111000010;
    16'b0010001000000001: out_v[318] = 10'b0110011000;
    16'b0000000000000011: out_v[318] = 10'b0110100011;
    16'b0010001000010010: out_v[318] = 10'b0000010011;
    16'b0010001000011011: out_v[318] = 10'b0100011000;
    16'b0010000000000010: out_v[318] = 10'b0010110100;
    16'b1000001000011011: out_v[318] = 10'b0100011111;
    16'b0100001000000100: out_v[318] = 10'b1111100011;
    16'b0110000000000010: out_v[318] = 10'b0110110111;
    16'b0100001000000000: out_v[318] = 10'b0111110000;
    16'b0110001000000010: out_v[318] = 10'b0110110011;
    16'b0010001000000110: out_v[318] = 10'b1011100010;
    16'b0100000000010011: out_v[318] = 10'b1100100101;
    16'b0110001000000100: out_v[318] = 10'b0011110111;
    16'b0001001000000010: out_v[318] = 10'b1100100001;
    16'b0001100000000010: out_v[318] = 10'b1011011011;
    16'b0001000000000000: out_v[318] = 10'b0011001100;
    16'b0000000000010110: out_v[318] = 10'b1101101100;
    16'b0001001000000000: out_v[318] = 10'b0110100110;
    16'b0000001000010110: out_v[318] = 10'b0111100101;
    16'b0001000000000010: out_v[318] = 10'b0001101011;
    16'b0001001000000100: out_v[318] = 10'b1101011010;
    16'b0010000000011001: out_v[318] = 10'b0100001110;
    16'b0000001000011001: out_v[318] = 10'b1101100111;
    16'b0010001000011001: out_v[318] = 10'b1111010011;
    16'b1010001000011001: out_v[318] = 10'b0011101101;
    16'b1010000000011001: out_v[318] = 10'b1011101101;
    16'b0000000000011001: out_v[318] = 10'b0110001110;
    16'b0010001000000101: out_v[318] = 10'b1011001011;
    16'b0010001000000111: out_v[318] = 10'b0110010010;
    16'b0100001000000010: out_v[318] = 10'b0111001110;
    default: out_v[318] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1100000010001110: out_v[319] = 10'b0010101101;
    16'b1100100010001110: out_v[319] = 10'b1000000111;
    16'b1100101010001110: out_v[319] = 10'b0110010011;
    16'b1000100010001010: out_v[319] = 10'b1011010010;
    16'b1100101010001100: out_v[319] = 10'b0110000101;
    16'b0100000010000110: out_v[319] = 10'b1011001001;
    16'b1000000000001010: out_v[319] = 10'b0000100001;
    16'b1000100010001110: out_v[319] = 10'b0001110011;
    16'b1100100010001010: out_v[319] = 10'b1000001111;
    16'b1100100000001010: out_v[319] = 10'b0110010101;
    16'b1000100000001010: out_v[319] = 10'b1110100110;
    16'b1000001000001000: out_v[319] = 10'b0101011011;
    16'b1100101000001100: out_v[319] = 10'b1100010111;
    16'b1100000010001100: out_v[319] = 10'b0010111100;
    16'b1100101000001000: out_v[319] = 10'b1001100011;
    16'b1000000010001110: out_v[319] = 10'b1011001111;
    16'b1100101010001000: out_v[319] = 10'b0001000011;
    16'b1100100000001000: out_v[319] = 10'b0011110110;
    16'b1100000000001100: out_v[319] = 10'b0100011011;
    16'b1100000000001010: out_v[319] = 10'b0010111100;
    16'b1000000010001100: out_v[319] = 10'b1100101110;
    16'b1100100000001110: out_v[319] = 10'b0001000111;
    16'b1100001010001100: out_v[319] = 10'b0111010011;
    16'b0100101010000100: out_v[319] = 10'b1011011110;
    16'b1100000000001110: out_v[319] = 10'b1011110000;
    16'b1100000010001010: out_v[319] = 10'b0100011011;
    16'b1000000000001000: out_v[319] = 10'b0001100101;
    16'b1000101010001100: out_v[319] = 10'b0011010011;
    16'b1000100000001000: out_v[319] = 10'b1001101110;
    16'b1100001000001000: out_v[319] = 10'b0101110110;
    16'b1000100000001110: out_v[319] = 10'b0110111011;
    16'b1000101000001000: out_v[319] = 10'b0100101101;
    16'b1100100010001100: out_v[319] = 10'b0000001110;
    16'b1000000010001010: out_v[319] = 10'b1111010000;
    16'b0100100010000110: out_v[319] = 10'b1111001010;
    16'b1000000000001110: out_v[319] = 10'b1001010111;
    16'b1100000000001000: out_v[319] = 10'b0011011110;
    16'b0000000000000100: out_v[319] = 10'b0101111010;
    16'b0000000000001100: out_v[319] = 10'b1101000111;
    16'b0000000010000100: out_v[319] = 10'b0011111110;
    16'b1100000000000000: out_v[319] = 10'b0111101110;
    16'b1000000000001100: out_v[319] = 10'b0101001101;
    16'b0000000010000000: out_v[319] = 10'b1101001001;
    16'b0100000000000000: out_v[319] = 10'b0111101111;
    16'b0000000000000000: out_v[319] = 10'b1010101100;
    16'b0000000010001100: out_v[319] = 10'b1011101110;
    16'b0000000000001000: out_v[319] = 10'b0100000010;
    16'b0000000000000010: out_v[319] = 10'b1001100100;
    16'b0100000000001000: out_v[319] = 10'b1001001101;
    16'b1100000010001000: out_v[319] = 10'b1101010110;
    16'b0100000000000010: out_v[319] = 10'b1001001010;
    16'b1000000010001000: out_v[319] = 10'b1000100101;
    16'b0100000010000000: out_v[319] = 10'b0000111111;
    16'b0100000010000100: out_v[319] = 10'b1010100111;
    16'b0100000000000100: out_v[319] = 10'b1111001001;
    16'b1000000000000000: out_v[319] = 10'b0000101010;
    16'b0000000010000110: out_v[319] = 10'b0110101101;
    16'b0000000000000110: out_v[319] = 10'b0001010101;
    16'b1101000000001100: out_v[319] = 10'b0111011001;
    16'b1001000000001000: out_v[319] = 10'b1101011011;
    16'b1101000000001000: out_v[319] = 10'b1111000101;
    16'b1101000000001010: out_v[319] = 10'b1101011110;
    16'b0000000010000010: out_v[319] = 10'b1000011100;
    16'b0000100000000010: out_v[319] = 10'b1110100000;
    16'b0000001000000010: out_v[319] = 10'b0100111010;
    16'b0100000010000010: out_v[319] = 10'b0011110010;
    16'b0100001000000010: out_v[319] = 10'b0100110100;
    16'b0000000000001010: out_v[319] = 10'b1010100001;
    16'b0000101000000010: out_v[319] = 10'b0011010110;
    16'b0100000010001110: out_v[319] = 10'b0110000011;
    16'b0100001000000000: out_v[319] = 10'b1001011011;
    16'b0100000010001010: out_v[319] = 10'b1100100111;
    16'b0000000010001010: out_v[319] = 10'b0001111010;
    16'b0000100010000010: out_v[319] = 10'b0001110010;
    16'b0100000000000110: out_v[319] = 10'b1001011010;
    16'b0000101000000000: out_v[319] = 10'b0011010010;
    16'b0100000000001010: out_v[319] = 10'b0100010101;
    16'b0000001000000000: out_v[319] = 10'b1111101011;
    16'b0000000010001110: out_v[319] = 10'b0100010001;
    16'b0100101000000010: out_v[319] = 10'b0101011001;
    16'b1100001010001110: out_v[319] = 10'b0001111000;
    16'b1000001000001010: out_v[319] = 10'b0111100000;
    16'b0000000010010110: out_v[319] = 10'b0111101011;
    16'b0000100010010010: out_v[319] = 10'b0011011011;
    16'b0000000010010010: out_v[319] = 10'b1011010010;
    16'b0000000010010100: out_v[319] = 10'b1100011011;
    16'b0000000000010100: out_v[319] = 10'b0010100010;
    16'b0000100010000110: out_v[319] = 10'b1010001000;
    16'b0000100000000000: out_v[319] = 10'b0101101111;
    16'b0000000000010010: out_v[319] = 10'b1101000100;
    16'b0000100010010110: out_v[319] = 10'b0001101000;
    16'b0000000000010110: out_v[319] = 10'b0111011101;
    16'b0100001010000100: out_v[319] = 10'b0110110110;
    16'b0100000010001100: out_v[319] = 10'b1100110101;
    16'b1000100010001100: out_v[319] = 10'b0110100110;
    16'b0000001010000100: out_v[319] = 10'b1010000100;
    16'b0000100010000100: out_v[319] = 10'b1100000111;
    16'b0100100010001100: out_v[319] = 10'b0101110100;
    16'b0100100010000100: out_v[319] = 10'b0100111010;
    16'b0000101010000100: out_v[319] = 10'b1110010111;
    16'b0100000000001100: out_v[319] = 10'b1110100010;
    16'b0000000010001000: out_v[319] = 10'b0100101101;
    16'b1000100010001000: out_v[319] = 10'b0100001010;
    16'b0100000010001000: out_v[319] = 10'b1110011011;
    16'b0000001010000110: out_v[319] = 10'b1001110011;
    16'b0100001010000110: out_v[319] = 10'b1000111010;
    16'b0100101010000110: out_v[319] = 10'b1110000101;
    default: out_v[319] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0110000000100000: out_v[320] = 10'b1011101111;
    16'b0010000000000001: out_v[320] = 10'b1000111111;
    16'b0100000101000001: out_v[320] = 10'b1110101101;
    16'b0000000000000001: out_v[320] = 10'b1001011010;
    16'b0100010000001000: out_v[320] = 10'b0001001111;
    16'b0101010100001001: out_v[320] = 10'b1010100100;
    16'b0010010000100001: out_v[320] = 10'b1010010101;
    16'b0100010000000000: out_v[320] = 10'b0011000101;
    16'b0010000001100001: out_v[320] = 10'b1101000101;
    16'b0110000000000001: out_v[320] = 10'b0111110101;
    16'b0111000100000001: out_v[320] = 10'b0110100111;
    16'b0101000100000001: out_v[320] = 10'b1001111001;
    16'b1111000100000001: out_v[320] = 10'b0011011111;
    16'b0100010000001001: out_v[320] = 10'b1011010010;
    16'b0000000000000000: out_v[320] = 10'b0111000001;
    16'b0100000100000001: out_v[320] = 10'b1111001010;
    16'b0110000000100001: out_v[320] = 10'b0011001110;
    16'b0101010100000001: out_v[320] = 10'b0011011111;
    16'b0100010000000001: out_v[320] = 10'b1011001111;
    16'b1101000100000001: out_v[320] = 10'b0101001101;
    16'b0100000000000000: out_v[320] = 10'b0111010001;
    16'b0111000100100001: out_v[320] = 10'b1101100001;
    16'b0100110000001000: out_v[320] = 10'b1001101010;
    16'b1101000000000001: out_v[320] = 10'b1001001011;
    16'b0110010000000001: out_v[320] = 10'b0010110001;
    16'b0110000001100001: out_v[320] = 10'b1100000101;
    16'b0100010100001001: out_v[320] = 10'b1111101000;
    16'b0000010000011000: out_v[320] = 10'b0011100011;
    16'b0100010000011000: out_v[320] = 10'b1011101001;
    16'b0000000100000001: out_v[320] = 10'b1001110011;
    16'b1101000100000000: out_v[320] = 10'b0111110000;
    16'b0010000000100001: out_v[320] = 10'b0111000111;
    16'b0100000000000001: out_v[320] = 10'b1101100011;
    16'b0110010000100001: out_v[320] = 10'b1011110111;
    16'b0100110000001001: out_v[320] = 10'b1000101110;
    16'b0101000000000001: out_v[320] = 10'b1000110111;
    16'b1111000100100001: out_v[320] = 10'b0101001011;
    16'b0100010100000001: out_v[320] = 10'b0111010110;
    16'b0100000100000000: out_v[320] = 10'b1101010100;
    16'b0101000100000000: out_v[320] = 10'b1000111000;
    16'b0110000100000001: out_v[320] = 10'b0011011000;
    16'b0010010001100001: out_v[320] = 10'b0110010011;
    16'b0010010001101001: out_v[320] = 10'b0011000011;
    16'b0100010000010000: out_v[320] = 10'b1101110011;
    16'b0010000001100000: out_v[320] = 10'b0011111000;
    16'b0000000001000000: out_v[320] = 10'b1100001110;
    16'b1100000001000000: out_v[320] = 10'b0101010001;
    16'b0101000001000000: out_v[320] = 10'b1001100110;
    16'b0100000001000000: out_v[320] = 10'b1100010100;
    16'b0101000000000000: out_v[320] = 10'b1101000111;
    16'b0001000001000000: out_v[320] = 10'b0011111110;
    16'b0000000001100000: out_v[320] = 10'b0001111011;
    16'b1101000001000000: out_v[320] = 10'b1001100110;
    16'b0100000001100000: out_v[320] = 10'b0000111111;
    16'b0010010001100000: out_v[320] = 10'b1010110010;
    16'b1101000000000000: out_v[320] = 10'b0101110100;
    16'b0000010001000000: out_v[320] = 10'b0101100110;
    16'b1000000001000000: out_v[320] = 10'b0001110111;
    16'b0100000101000000: out_v[320] = 10'b0100100011;
    16'b0101000001100000: out_v[320] = 10'b1010011001;
    16'b0110000100100001: out_v[320] = 10'b0001010110;
    16'b0110000101100001: out_v[320] = 10'b1001110100;
    16'b0110000000000000: out_v[320] = 10'b1001010100;
    16'b0000000100000000: out_v[320] = 10'b0000011111;
    16'b0010000100100001: out_v[320] = 10'b1111000110;
    16'b0010000000100000: out_v[320] = 10'b1001101010;
    16'b0110000100110001: out_v[320] = 10'b1110010101;
    16'b0110010100110000: out_v[320] = 10'b1101110101;
    16'b0111000101100001: out_v[320] = 10'b1110100011;
    16'b0010000101100001: out_v[320] = 10'b0101011000;
    16'b0110000101100000: out_v[320] = 10'b1000010011;
    16'b0110010000110001: out_v[320] = 10'b1011110111;
    16'b0110000100100000: out_v[320] = 10'b1011001001;
    16'b0110000000110001: out_v[320] = 10'b1111010011;
    16'b0000000101000000: out_v[320] = 10'b0110010111;
    16'b0110010100100001: out_v[320] = 10'b1011101010;
    16'b0110010100110001: out_v[320] = 10'b1100100111;
    16'b0110000001100000: out_v[320] = 10'b0111010110;
    16'b0111000101100000: out_v[320] = 10'b1101001010;
    16'b0110010000110000: out_v[320] = 10'b1111010010;
    16'b0101000101000000: out_v[320] = 10'b0111001101;
    16'b1101000101000000: out_v[320] = 10'b1101001001;
    16'b1111000000100000: out_v[320] = 10'b0110010011;
    16'b1111000101100000: out_v[320] = 10'b0010001100;
    16'b1101000101100000: out_v[320] = 10'b1101010110;
    16'b0100010001100000: out_v[320] = 10'b0000011111;
    16'b1101000001100000: out_v[320] = 10'b1001001111;
    16'b1111000001100000: out_v[320] = 10'b1011100111;
    16'b1101000100100000: out_v[320] = 10'b0110011010;
    16'b0100000001010000: out_v[320] = 10'b1011110000;
    16'b1111000100100000: out_v[320] = 10'b0010110001;
    16'b0110010001100000: out_v[320] = 10'b0000011011;
    16'b0100000000100000: out_v[320] = 10'b1101110001;
    16'b1101000000100000: out_v[320] = 10'b0101011000;
    16'b0100010001110000: out_v[320] = 10'b1111100110;
    16'b0100000001100001: out_v[320] = 10'b1011011111;
    16'b0101000101100000: out_v[320] = 10'b1111011011;
    16'b0100000001000001: out_v[320] = 10'b0011111001;
    16'b0100010001000000: out_v[320] = 10'b1011110100;
    16'b0101000101010000: out_v[320] = 10'b1100011111;
    16'b0100000101100000: out_v[320] = 10'b1110110101;
    16'b0101000101000001: out_v[320] = 10'b1011001010;
    16'b0100010001010000: out_v[320] = 10'b1101010110;
    16'b0011000000100000: out_v[320] = 10'b1011101101;
    16'b0000000000100000: out_v[320] = 10'b1101001000;
    16'b0010000100100000: out_v[320] = 10'b0011011101;
    16'b0110010000100000: out_v[320] = 10'b1011101011;
    16'b1011010000100000: out_v[320] = 10'b1111011011;
    16'b0001000000100000: out_v[320] = 10'b0100010010;
    16'b0010010000101000: out_v[320] = 10'b1100010011;
    16'b0111000000100000: out_v[320] = 10'b1010110001;
    16'b1110000000100000: out_v[320] = 10'b1101101000;
    16'b1001000001100000: out_v[320] = 10'b1100010100;
    16'b0010010000100000: out_v[320] = 10'b0010100100;
    16'b1011000000100000: out_v[320] = 10'b0011100011;
    16'b0011000001100000: out_v[320] = 10'b1011011011;
    16'b1001000000100000: out_v[320] = 10'b0011110110;
    16'b0010000000101000: out_v[320] = 10'b1010011010;
    16'b0010000101100000: out_v[320] = 10'b1001000101;
    16'b0010100000101000: out_v[320] = 10'b0000111111;
    16'b1010000000100000: out_v[320] = 10'b1111011100;
    16'b0011000000100001: out_v[320] = 10'b0101111010;
    16'b1011000001100000: out_v[320] = 10'b0110110000;
    16'b1010000001100000: out_v[320] = 10'b1011011101;
    16'b1010010000100000: out_v[320] = 10'b0101001110;
    16'b0110000000101000: out_v[320] = 10'b0011111111;
    16'b0000010000100000: out_v[320] = 10'b0001011100;
    16'b1111010000100000: out_v[320] = 10'b0000111100;
    16'b0110010000101000: out_v[320] = 10'b0111100111;
    16'b0010000000000000: out_v[320] = 10'b1101101000;
    16'b1111010100100000: out_v[320] = 10'b0110110111;
    16'b0111000100100000: out_v[320] = 10'b0011110011;
    16'b0000010000101000: out_v[320] = 10'b1001001011;
    16'b0010010001101000: out_v[320] = 10'b0000110100;
    16'b0000100001101000: out_v[320] = 10'b0011010001;
    16'b0000100000101000: out_v[320] = 10'b1101101100;
    16'b0000100001001001: out_v[320] = 10'b0001110111;
    16'b0101000000100000: out_v[320] = 10'b0010110011;
    16'b0000010000001000: out_v[320] = 10'b0111101100;
    16'b0000010000000000: out_v[320] = 10'b0111010011;
    16'b0101000100100000: out_v[320] = 10'b0110110001;
    16'b0010100001101000: out_v[320] = 10'b0111110001;
    16'b0000100001101001: out_v[320] = 10'b1011101110;
    16'b0010000100000001: out_v[320] = 10'b1101011010;
    16'b0110000100000000: out_v[320] = 10'b1000101001;
    16'b0010000100000000: out_v[320] = 10'b1001001111;
    16'b1001000101000000: out_v[320] = 10'b1010011111;
    16'b1001000000000000: out_v[320] = 10'b0111111100;
    16'b1000000000000000: out_v[320] = 10'b0110111101;
    16'b1001000001000000: out_v[320] = 10'b0010110110;
    16'b0000010001001000: out_v[320] = 10'b0011000111;
    16'b0000000010000000: out_v[320] = 10'b0101110110;
    16'b0000000000001000: out_v[320] = 10'b0111101100;
    16'b0000010010001000: out_v[320] = 10'b0110010111;
    16'b1001001000000000: out_v[320] = 10'b1111111111;
    16'b0000001000000000: out_v[320] = 10'b1111110111;
    16'b1100000000000000: out_v[320] = 10'b0001110110;
    16'b1000001000000000: out_v[320] = 10'b1110110101;
    16'b1001001001000000: out_v[320] = 10'b0101010101;
    16'b0000000001001000: out_v[320] = 10'b1010000100;
    16'b0110100000101001: out_v[320] = 10'b1110101111;
    16'b1111000000100001: out_v[320] = 10'b0111010011;
    16'b1111010001100000: out_v[320] = 10'b1011100110;
    16'b0111000001100001: out_v[320] = 10'b1110010100;
    16'b1101010000100000: out_v[320] = 10'b0011010111;
    16'b1111010000100001: out_v[320] = 10'b0110110001;
    16'b1111000101100001: out_v[320] = 10'b0001100011;
    16'b0100010000100000: out_v[320] = 10'b1000011011;
    16'b0010100000101001: out_v[320] = 10'b1110100001;
    16'b0110100001101001: out_v[320] = 10'b1100011010;
    16'b0110110000101001: out_v[320] = 10'b1010100011;
    16'b1111000001100001: out_v[320] = 10'b1111100111;
    16'b0110010000101001: out_v[320] = 10'b0000110110;
    16'b0010010000101001: out_v[320] = 10'b0011101110;
    16'b0010110000101001: out_v[320] = 10'b0111011010;
    16'b0110010001101001: out_v[320] = 10'b1110000111;
    16'b0110010001100001: out_v[320] = 10'b0100100000;
    16'b0111000001100000: out_v[320] = 10'b0111010000;
    16'b1100000001100000: out_v[320] = 10'b1011100011;
    16'b1000000000100000: out_v[320] = 10'b1100100011;
    16'b0111000000000000: out_v[320] = 10'b1101001001;
    16'b1000000001100000: out_v[320] = 10'b1001100111;
    16'b1100000000100000: out_v[320] = 10'b1100100111;
    16'b1111000000000000: out_v[320] = 10'b1001101011;
    16'b1110000001100000: out_v[320] = 10'b0011000010;
    default: out_v[320] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001010000100001: out_v[321] = 10'b1010001011;
    16'b0001000000100001: out_v[321] = 10'b0011011100;
    16'b0001000001100001: out_v[321] = 10'b0110110101;
    16'b0000000000100001: out_v[321] = 10'b1000000101;
    16'b0001000001000001: out_v[321] = 10'b1011011001;
    16'b0000000000000001: out_v[321] = 10'b1000101011;
    16'b0001000001000000: out_v[321] = 10'b1100100110;
    16'b0001000000000001: out_v[321] = 10'b0011010011;
    16'b0000010000100001: out_v[321] = 10'b0010100101;
    16'b0000000001100001: out_v[321] = 10'b0110101001;
    16'b0000000000000000: out_v[321] = 10'b1100000101;
    16'b0000000000100000: out_v[321] = 10'b1010101001;
    16'b0001000001100000: out_v[321] = 10'b1011100110;
    16'b0001000000000000: out_v[321] = 10'b1100110101;
    16'b0001000001100101: out_v[321] = 10'b0011100110;
    16'b0000010000000001: out_v[321] = 10'b0011100001;
    16'b0001010000000001: out_v[321] = 10'b1000100111;
    16'b0001000000100000: out_v[321] = 10'b1101000110;
    16'b0001010001100001: out_v[321] = 10'b1000111010;
    16'b0000010000100000: out_v[321] = 10'b1101001011;
    16'b0000010000000000: out_v[321] = 10'b1001101101;
    16'b0000000001100000: out_v[321] = 10'b0101011101;
    16'b0001010000100000: out_v[321] = 10'b0001011111;
    16'b0000000001000100: out_v[321] = 10'b0010100010;
    16'b0000000000000100: out_v[321] = 10'b0110000011;
    16'b0000010001000100: out_v[321] = 10'b0011010111;
    16'b0001000001000100: out_v[321] = 10'b1001100110;
    16'b0000000001100100: out_v[321] = 10'b1100011011;
    16'b0000000001000101: out_v[321] = 10'b0111011010;
    16'b0000000001000000: out_v[321] = 10'b1001101100;
    16'b0000000000100100: out_v[321] = 10'b1111011011;
    16'b0000000001001100: out_v[321] = 10'b1011100100;
    16'b0001000001101100: out_v[321] = 10'b0011110011;
    16'b0001000000000100: out_v[321] = 10'b0010101001;
    16'b0001000001001100: out_v[321] = 10'b1111100101;
    16'b0001000001100100: out_v[321] = 10'b0111001100;
    16'b0000000000001110: out_v[321] = 10'b0001110110;
    16'b0001000001001000: out_v[321] = 10'b1100101110;
    16'b0000000001001110: out_v[321] = 10'b1101101011;
    16'b0000000001001000: out_v[321] = 10'b0111010000;
    16'b0000000000001100: out_v[321] = 10'b1010100010;
    16'b0001000000100100: out_v[321] = 10'b1110011010;
    16'b0001000001101000: out_v[321] = 10'b1101011110;
    16'b0000000001001010: out_v[321] = 10'b1100100101;
    16'b0001000001001110: out_v[321] = 10'b1101111111;
    16'b0001000001001010: out_v[321] = 10'b0100001010;
    16'b0000000001000001: out_v[321] = 10'b1100101101;
    16'b0001000001000101: out_v[321] = 10'b0110010010;
    16'b0001010000000000: out_v[321] = 10'b0110010011;
    16'b0001000000000101: out_v[321] = 10'b0001111100;
    16'b0001010000000100: out_v[321] = 10'b0001111010;
    16'b0000010000100100: out_v[321] = 10'b0001001100;
    16'b0001010000000101: out_v[321] = 10'b1100100110;
    16'b0001000000100101: out_v[321] = 10'b0100001110;
    16'b0000010000000100: out_v[321] = 10'b0101001100;
    16'b0000010000000101: out_v[321] = 10'b0101000110;
    16'b0000000000000101: out_v[321] = 10'b0001010101;
    16'b0001010000100101: out_v[321] = 10'b1101000100;
    16'b0001010000100100: out_v[321] = 10'b1100001010;
    16'b0000010001100101: out_v[321] = 10'b1000111011;
    16'b0000010001000101: out_v[321] = 10'b0001111001;
    16'b0000010001000001: out_v[321] = 10'b0110001100;
    16'b0000000001100101: out_v[321] = 10'b1001010000;
    16'b0001010001100101: out_v[321] = 10'b1100100110;
    16'b0000000000100101: out_v[321] = 10'b1100010010;
    16'b0001010001000101: out_v[321] = 10'b1100010000;
    16'b0011000000100000: out_v[321] = 10'b1100100000;
    16'b0001010001000001: out_v[321] = 10'b0110011000;
    16'b0000010001100001: out_v[321] = 10'b0110101000;
    16'b0001001001000101: out_v[321] = 10'b0110011111;
    16'b0001001001000001: out_v[321] = 10'b1100110111;
    16'b0001001001000000: out_v[321] = 10'b1101111010;
    16'b0001001001000100: out_v[321] = 10'b0100101111;
    16'b0000010001000000: out_v[321] = 10'b1111010010;
    16'b0011000000100001: out_v[321] = 10'b1110100111;
    16'b1000010001100000: out_v[321] = 10'b1111011010;
    16'b0011000000000000: out_v[321] = 10'b1110100011;
    16'b1000010001000001: out_v[321] = 10'b0111111110;
    16'b1000010001100001: out_v[321] = 10'b0111010001;
    16'b0001010001100000: out_v[321] = 10'b0110110010;
    16'b0010000000000000: out_v[321] = 10'b1111001010;
    16'b1000010001000000: out_v[321] = 10'b1101110011;
    16'b1000010000000000: out_v[321] = 10'b1100101111;
    16'b0000010001100000: out_v[321] = 10'b0100001110;
    16'b1000010000000001: out_v[321] = 10'b0111111011;
    16'b1011010000100000: out_v[321] = 10'b1111011111;
    16'b1001010001100001: out_v[321] = 10'b0111101111;
    16'b0001010001000100: out_v[321] = 10'b0010101000;
    16'b1001010000100001: out_v[321] = 10'b0110001111;
    16'b0011010000100000: out_v[321] = 10'b1111100011;
    16'b1011010001100000: out_v[321] = 10'b1101111011;
    16'b0011000000000001: out_v[321] = 10'b0111011010;
    16'b1001010000100000: out_v[321] = 10'b1111110100;
    16'b0001010001000000: out_v[321] = 10'b0010010001;
    16'b1000010001000100: out_v[321] = 10'b1011100101;
    16'b1001010001100000: out_v[321] = 10'b1001111101;
    16'b0000010000100101: out_v[321] = 10'b0111000100;
    16'b0000010001100100: out_v[321] = 10'b0111110001;
    16'b1000010001100101: out_v[321] = 10'b1000001100;
    16'b1000010000100101: out_v[321] = 10'b1101111110;
    16'b1001010000100101: out_v[321] = 10'b1101010111;
    16'b1000010001000101: out_v[321] = 10'b1101101111;
    default: out_v[321] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010010110101110: out_v[322] = 10'b1010101111;
    16'b0001010110101110: out_v[322] = 10'b0110111101;
    16'b0001010110101010: out_v[322] = 10'b0000110111;
    16'b0011010100101010: out_v[322] = 10'b0011101011;
    16'b0011010100101110: out_v[322] = 10'b1011110001;
    16'b0000010110101110: out_v[322] = 10'b1010110111;
    16'b0010000110101000: out_v[322] = 10'b0010100011;
    16'b0011000110101000: out_v[322] = 10'b0110010100;
    16'b0011010110101110: out_v[322] = 10'b0101101011;
    16'b0011010000101010: out_v[322] = 10'b0010010111;
    16'b0011010100001110: out_v[322] = 10'b0111100011;
    16'b0011000100101100: out_v[322] = 10'b1101011110;
    16'b0001000110101010: out_v[322] = 10'b1101001000;
    16'b0011010110100110: out_v[322] = 10'b1011000111;
    16'b0011010110101010: out_v[322] = 10'b0111000100;
    16'b0010000100101000: out_v[322] = 10'b1001010111;
    16'b0011010010101010: out_v[322] = 10'b1011101011;
    16'b0011010100001010: out_v[322] = 10'b0010100011;
    16'b0010010110111110: out_v[322] = 10'b1010000111;
    16'b0010010100001110: out_v[322] = 10'b1000010101;
    16'b0001000110101000: out_v[322] = 10'b1111100110;
    16'b0011000100101000: out_v[322] = 10'b1110010111;
    16'b0011010000001110: out_v[322] = 10'b1000111110;
    16'b0001000110101100: out_v[322] = 10'b1001011111;
    16'b0000000110101000: out_v[322] = 10'b1010000101;
    16'b0011000000001000: out_v[322] = 10'b0000001011;
    16'b0011000000001010: out_v[322] = 10'b1110111110;
    16'b0011000110101100: out_v[322] = 10'b1110001001;
    16'b0001000110101110: out_v[322] = 10'b0001111111;
    16'b0011000110101010: out_v[322] = 10'b0100011110;
    16'b0010010100101110: out_v[322] = 10'b1000010111;
    16'b0011000100001000: out_v[322] = 10'b1110111011;
    16'b0011010000001010: out_v[322] = 10'b0111100110;
    16'b0011010110111110: out_v[322] = 10'b1110100011;
    16'b0001010110111110: out_v[322] = 10'b0010011110;
    16'b0011010010101110: out_v[322] = 10'b0001111011;
    16'b0011000000101010: out_v[322] = 10'b1110111100;
    16'b0011000100101010: out_v[322] = 10'b0110100110;
    16'b0011000000101000: out_v[322] = 10'b1010011111;
    16'b0011010000101110: out_v[322] = 10'b0011110101;
    16'b0011000110101110: out_v[322] = 10'b1111110110;
    16'b0000010000011010: out_v[322] = 10'b1000100011;
    16'b0010000010100000: out_v[322] = 10'b0010110111;
    16'b0010000010010000: out_v[322] = 10'b1101011001;
    16'b0000000000011000: out_v[322] = 10'b1011110011;
    16'b0010000010111000: out_v[322] = 10'b1010100011;
    16'b0010000010110000: out_v[322] = 10'b1000111110;
    16'b0010000110100000: out_v[322] = 10'b0101010011;
    16'b0000000010010000: out_v[322] = 10'b1001011100;
    16'b0000000000011010: out_v[322] = 10'b1101110001;
    16'b0010000000011000: out_v[322] = 10'b1010100100;
    16'b0000000010110000: out_v[322] = 10'b1110000101;
    16'b0000000010100000: out_v[322] = 10'b0000001111;
    16'b0000010010011010: out_v[322] = 10'b1000100110;
    16'b0010000110110000: out_v[322] = 10'b0011110011;
    16'b0000000010011000: out_v[322] = 10'b0001110100;
    16'b0000000000010000: out_v[322] = 10'b0000110010;
    16'b0000000010111000: out_v[322] = 10'b0111111101;
    16'b0000010000010010: out_v[322] = 10'b0001110011;
    16'b0010000010011000: out_v[322] = 10'b1101100011;
    16'b0000000000001000: out_v[322] = 10'b1101101011;
    16'b0000000000000000: out_v[322] = 10'b0001010111;
    16'b0000000000010010: out_v[322] = 10'b0001111001;
    16'b0010000010000000: out_v[322] = 10'b1110011101;
    16'b0000000010011010: out_v[322] = 10'b0000110111;
    16'b0010000000000000: out_v[322] = 10'b1110100011;
    16'b0000000110100000: out_v[322] = 10'b1001010111;
    16'b0010000110111000: out_v[322] = 10'b0010010110;
    16'b0010000000001000: out_v[322] = 10'b0111000101;
    16'b0010000010101000: out_v[322] = 10'b1110011011;
    16'b0010010100011110: out_v[322] = 10'b1100100111;
    16'b0010000100001000: out_v[322] = 10'b1000100011;
    16'b0010000100011010: out_v[322] = 10'b1101100011;
    16'b0010010100111010: out_v[322] = 10'b0010011101;
    16'b0010010100011010: out_v[322] = 10'b0111101101;
    16'b0010000100011000: out_v[322] = 10'b1100110101;
    16'b0010010000001010: out_v[322] = 10'b0001001101;
    16'b0000000000110000: out_v[322] = 10'b1001100001;
    16'b0010010100010110: out_v[322] = 10'b1111000110;
    16'b0010000000011010: out_v[322] = 10'b1111010100;
    16'b0010000000010000: out_v[322] = 10'b1011111101;
    16'b0010010100111110: out_v[322] = 10'b1111111110;
    16'b0011010100011110: out_v[322] = 10'b1011110111;
    16'b0010010100110010: out_v[322] = 10'b0111111111;
    16'b0011010100111110: out_v[322] = 10'b0010011111;
    16'b0010000100010000: out_v[322] = 10'b1000100111;
    16'b0010010100001010: out_v[322] = 10'b1100011100;
    16'b0010010000011110: out_v[322] = 10'b0110001001;
    16'b0010010000001110: out_v[322] = 10'b1010011011;
    16'b0010000100111000: out_v[322] = 10'b1011111101;
    16'b0010010100101010: out_v[322] = 10'b0011011101;
    16'b0010010000111110: out_v[322] = 10'b1101001010;
    16'b0011010100010110: out_v[322] = 10'b1011100000;
    16'b0000000110110000: out_v[322] = 10'b0001011110;
    16'b0010010000011010: out_v[322] = 10'b0110000010;
    16'b1010000100011000: out_v[322] = 10'b1110011001;
    16'b0010010000111010: out_v[322] = 10'b0100010000;
    16'b0010010000101010: out_v[322] = 10'b1000110111;
    16'b0010010100010010: out_v[322] = 10'b0100000111;
    16'b0010010110111010: out_v[322] = 10'b1110000100;
    16'b0011010000011110: out_v[322] = 10'b1001011101;
    16'b0010000110011000: out_v[322] = 10'b0110011111;
    16'b0011010000111110: out_v[322] = 10'b0111110011;
    16'b0010000110000100: out_v[322] = 10'b0111111001;
    16'b0010010110001110: out_v[322] = 10'b1011001010;
    16'b0010000110111100: out_v[322] = 10'b1001101010;
    16'b0010000110011100: out_v[322] = 10'b1111011011;
    16'b0010000110101100: out_v[322] = 10'b1111111000;
    16'b0010000010001100: out_v[322] = 10'b1001100111;
    16'b0010000000011100: out_v[322] = 10'b1011101110;
    16'b0010000110001100: out_v[322] = 10'b1110010001;
    16'b0010000100011100: out_v[322] = 10'b0010101011;
    16'b0010000000000100: out_v[322] = 10'b1101110100;
    16'b0010000100000000: out_v[322] = 10'b0101100100;
    16'b0010010110001100: out_v[322] = 10'b1110111110;
    16'b0010000110000000: out_v[322] = 10'b1000001101;
    16'b0010000010101100: out_v[322] = 10'b0111011001;
    16'b0010000110010000: out_v[322] = 10'b1111001101;
    16'b0010000110001110: out_v[322] = 10'b1001001111;
    16'b0000000100110000: out_v[322] = 10'b1101101101;
    16'b0010000100001100: out_v[322] = 10'b0001110100;
    16'b0010000010000100: out_v[322] = 10'b1111010111;
    16'b0010000110001000: out_v[322] = 10'b1011001100;
    16'b0010000100001010: out_v[322] = 10'b1110001011;
    16'b0010000000001100: out_v[322] = 10'b1011111010;
    16'b0000010100010110: out_v[322] = 10'b0000011110;
    16'b0000000100010100: out_v[322] = 10'b0101010011;
    16'b0000000100010000: out_v[322] = 10'b0001010011;
    16'b0001010010111110: out_v[322] = 10'b1001101101;
    16'b0000010000011110: out_v[322] = 10'b1000010101;
    16'b0000010010110010: out_v[322] = 10'b1001011001;
    16'b0000000110110100: out_v[322] = 10'b0011001011;
    16'b0000010100010010: out_v[322] = 10'b0010100101;
    16'b0010000110110100: out_v[322] = 10'b0011101000;
    16'b0001010000011110: out_v[322] = 10'b1011111110;
    16'b0001010100000110: out_v[322] = 10'b1011001011;
    16'b0000010100000010: out_v[322] = 10'b0110110011;
    16'b0000000100000000: out_v[322] = 10'b0001011011;
    16'b0000010000010110: out_v[322] = 10'b0111011000;
    16'b0000010100000110: out_v[322] = 10'b0111010000;
    16'b0001010100010110: out_v[322] = 10'b0000111101;
    16'b0000010000000010: out_v[322] = 10'b0100110010;
    16'b0000010010111010: out_v[322] = 10'b1101011101;
    16'b0000010100110110: out_v[322] = 10'b0101100001;
    16'b0001010110110110: out_v[322] = 10'b1001011111;
    16'b0001010000010110: out_v[322] = 10'b0010011010;
    16'b0001010100110110: out_v[322] = 10'b0000111111;
    16'b0000010000110110: out_v[322] = 10'b1001000110;
    16'b0000010010111110: out_v[322] = 10'b0010110111;
    16'b0000010110110110: out_v[322] = 10'b1010010010;
    16'b0000010010110110: out_v[322] = 10'b1001111010;
    16'b0000000000010100: out_v[322] = 10'b0000111111;
    16'b0000000010110100: out_v[322] = 10'b0010111001;
    16'b0000010000000110: out_v[322] = 10'b1101011011;
    16'b0000000000010110: out_v[322] = 10'b0111101000;
    16'b0010010110110110: out_v[322] = 10'b0010010011;
    16'b0000010010011110: out_v[322] = 10'b1100010011;
    16'b0001010010011010: out_v[322] = 10'b1101110000;
    16'b0000000010101000: out_v[322] = 10'b0001111110;
    16'b0000000110111010: out_v[322] = 10'b1011110010;
    16'b0000000100111000: out_v[322] = 10'b0110010110;
    16'b0000000110101100: out_v[322] = 10'b0001110000;
    16'b0000000100101100: out_v[322] = 10'b0010101010;
    16'b0000000110111000: out_v[322] = 10'b1010111101;
    16'b0000000000100100: out_v[322] = 10'b1101111111;
    16'b0010000000111100: out_v[322] = 10'b1011010010;
    16'b0010000100110000: out_v[322] = 10'b0110101100;
    16'b0000000110111100: out_v[322] = 10'b0001011110;
    16'b0000000010111010: out_v[322] = 10'b0111100000;
    16'b0010000100111100: out_v[322] = 10'b1011111000;
    16'b0010000100100000: out_v[322] = 10'b0011111010;
    16'b0000000110011000: out_v[322] = 10'b1101000011;
    16'b0000000100100000: out_v[322] = 10'b0110100101;
    16'b0000000010001010: out_v[322] = 10'b1100011110;
    16'b0010000100101100: out_v[322] = 10'b0111110000;
    16'b0010000000101100: out_v[322] = 10'b0001110000;
    16'b0100000101110000: out_v[322] = 10'b1001110111;
    16'b0000000100101000: out_v[322] = 10'b0110110011;
    16'b0100000111110000: out_v[322] = 10'b0010001111;
    16'b0000000100000100: out_v[322] = 10'b1101101011;
    16'b0010010100101100: out_v[322] = 10'b0100000111;
    16'b0010000100010100: out_v[322] = 10'b0111110001;
    16'b0000010110111100: out_v[322] = 10'b0011000101;
    16'b0010010110111100: out_v[322] = 10'b1010111001;
    16'b0000000110011100: out_v[322] = 10'b1001000010;
    16'b0010000100100100: out_v[322] = 10'b1101001111;
    16'b0001010100000010: out_v[322] = 10'b1101101011;
    16'b0010010110101100: out_v[322] = 10'b0111011000;
    16'b0001010100011010: out_v[322] = 10'b1011111111;
    16'b0001010100001010: out_v[322] = 10'b1101100010;
    16'b0010000110100100: out_v[322] = 10'b1111001110;
    16'b0010000100110100: out_v[322] = 10'b0111101011;
    16'b0010010100111100: out_v[322] = 10'b0010110011;
    16'b0010000100000100: out_v[322] = 10'b1101100101;
    16'b0001010110000110: out_v[322] = 10'b0111001100;
    16'b0101010010101110: out_v[322] = 10'b0111111110;
    16'b0001010110100110: out_v[322] = 10'b1110001110;
    16'b0100010011101110: out_v[322] = 10'b0110011011;
    16'b0100010001101010: out_v[322] = 10'b0111101011;
    16'b0000010100100110: out_v[322] = 10'b0010001000;
    16'b0000010110100010: out_v[322] = 10'b0011001011;
    16'b0100010111100110: out_v[322] = 10'b1001010011;
    16'b0000010110100110: out_v[322] = 10'b0011010110;
    16'b0100010111101110: out_v[322] = 10'b1111010011;
    16'b0000010100100010: out_v[322] = 10'b1011010000;
    16'b0100010011100010: out_v[322] = 10'b0111010100;
    16'b0100010001100010: out_v[322] = 10'b1101101101;
    16'b0101010011101110: out_v[322] = 10'b0100111111;
    16'b0000010110000110: out_v[322] = 10'b0010000111;
    16'b0001010010101110: out_v[322] = 10'b0111000111;
    16'b0000010000101110: out_v[322] = 10'b1100111010;
    16'b0000010000101010: out_v[322] = 10'b0001010111;
    16'b0000000000100000: out_v[322] = 10'b0111110100;
    16'b0100010110100110: out_v[322] = 10'b1110110011;
    16'b0101010111100110: out_v[322] = 10'b0111010010;
    16'b0100010011101010: out_v[322] = 10'b0001010110;
    16'b0000010010101010: out_v[322] = 10'b0011100001;
    16'b0100010000101010: out_v[322] = 10'b1111110011;
    16'b0100010011100110: out_v[322] = 10'b1111011010;
    16'b0000010000100010: out_v[322] = 10'b1011011111;
    16'b0101010011100110: out_v[322] = 10'b0101111111;
    16'b0101010111101110: out_v[322] = 10'b0010111100;
    16'b0000010010100010: out_v[322] = 10'b0111110111;
    16'b0000010010100110: out_v[322] = 10'b1111000111;
    16'b0100010001101110: out_v[322] = 10'b1101111101;
    16'b0001010000101110: out_v[322] = 10'b0010100010;
    16'b0101010110100110: out_v[322] = 10'b0110101100;
    16'b0001010010001110: out_v[322] = 10'b0111001101;
    16'b0100000001100000: out_v[322] = 10'b0110011011;
    16'b0100010010101010: out_v[322] = 10'b0000001101;
    16'b0000010010101110: out_v[322] = 10'b1001011010;
    16'b0101010001101110: out_v[322] = 10'b0011100011;
    16'b0100010001100110: out_v[322] = 10'b0101111111;
    16'b0100000001101000: out_v[322] = 10'b0111110001;
    16'b0000000000110100: out_v[322] = 10'b0110000011;
    16'b0100010101100110: out_v[322] = 10'b0111110101;
    16'b0011010100011010: out_v[322] = 10'b0110000000;
    16'b0011010110111010: out_v[322] = 10'b0101100010;
    16'b0000010110111010: out_v[322] = 10'b0110001101;
    16'b0010010010110010: out_v[322] = 10'b0101010001;
    16'b0010010010111010: out_v[322] = 10'b0000011111;
    16'b0000010100110010: out_v[322] = 10'b1110000011;
    16'b0010000110111010: out_v[322] = 10'b0011110100;
    16'b0000010100111010: out_v[322] = 10'b0101011110;
    16'b0001010010111010: out_v[322] = 10'b1111101100;
    16'b0011010010111110: out_v[322] = 10'b0111000100;
    16'b0001010010110010: out_v[322] = 10'b0010111111;
    16'b0000010000110010: out_v[322] = 10'b1101001011;
    16'b0010010110110010: out_v[322] = 10'b0111110110;
    16'b0000010000111010: out_v[322] = 10'b0111110011;
    16'b0010010110011010: out_v[322] = 10'b0011011111;
    16'b0011010010111010: out_v[322] = 10'b1001001001;
    16'b0010000100111010: out_v[322] = 10'b1010111111;
    16'b0011010100111010: out_v[322] = 10'b1011010100;
    16'b0011010010110010: out_v[322] = 10'b1011111000;
    16'b0010010000110010: out_v[322] = 10'b0110110110;
    16'b0100010011111110: out_v[322] = 10'b0011010110;
    16'b0100010000110010: out_v[322] = 10'b1000101111;
    16'b0100010011110010: out_v[322] = 10'b1101001010;
    16'b0101010111110110: out_v[322] = 10'b0111001111;
    16'b0000010000100110: out_v[322] = 10'b1001000110;
    16'b0100010011111010: out_v[322] = 10'b0101011111;
    16'b0100010011110110: out_v[322] = 10'b0001111011;
    16'b0101010011111110: out_v[322] = 10'b0101111110;
    16'b0000010110110010: out_v[322] = 10'b1111000101;
    16'b0100010001110010: out_v[322] = 10'b1001111111;
    16'b0100010001110110: out_v[322] = 10'b0111101110;
    16'b0000010100110100: out_v[322] = 10'b1001101111;
    16'b0000000100110100: out_v[322] = 10'b1011010101;
    16'b0101010001111110: out_v[322] = 10'b1001100111;
    16'b0101010011110110: out_v[322] = 10'b1000101111;
    16'b0001010100100110: out_v[322] = 10'b0101111010;
    16'b0100010001111010: out_v[322] = 10'b1111100011;
    default: out_v[322] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0101000000000011: out_v[323] = 10'b1101001001;
    16'b0111000000000011: out_v[323] = 10'b1000100100;
    16'b1111000000000011: out_v[323] = 10'b1010011110;
    16'b0111000000000000: out_v[323] = 10'b0100111101;
    16'b0111000000000001: out_v[323] = 10'b1001100001;
    16'b0110000000000001: out_v[323] = 10'b1111010000;
    16'b1111000000000001: out_v[323] = 10'b0010010001;
    16'b0100000000000001: out_v[323] = 10'b1011101110;
    16'b0111000000000010: out_v[323] = 10'b1001110010;
    16'b0011000000000111: out_v[323] = 10'b1110000100;
    16'b0111000000000111: out_v[323] = 10'b0000101111;
    16'b0110000000000111: out_v[323] = 10'b1111000001;
    16'b0110000000000010: out_v[323] = 10'b1000100111;
    16'b0011000000000001: out_v[323] = 10'b0110110100;
    16'b1011000000000010: out_v[323] = 10'b1001010110;
    16'b0110000000000011: out_v[323] = 10'b0110001111;
    16'b0111000100000011: out_v[323] = 10'b1001110101;
    16'b0010000000000001: out_v[323] = 10'b1001010111;
    16'b0101000000000001: out_v[323] = 10'b1101101001;
    16'b0011000000000010: out_v[323] = 10'b1011111100;
    16'b0011000000000011: out_v[323] = 10'b0010110100;
    16'b0101000000000010: out_v[323] = 10'b1100000011;
    16'b0011000000000000: out_v[323] = 10'b1011001110;
    16'b0110000000000000: out_v[323] = 10'b1101110000;
    16'b0001000000000010: out_v[323] = 10'b0111001110;
    16'b0111000100000111: out_v[323] = 10'b0111011111;
    16'b1111000000000111: out_v[323] = 10'b1100111011;
    16'b0010000000000011: out_v[323] = 10'b1000001111;
    16'b0001000000000110: out_v[323] = 10'b0101101110;
    16'b0000000000000010: out_v[323] = 10'b0111011000;
    16'b0001000000000000: out_v[323] = 10'b0001001111;
    16'b0010000000000000: out_v[323] = 10'b1111000000;
    16'b0001000000000100: out_v[323] = 10'b0111100110;
    16'b0000000000000011: out_v[323] = 10'b0111011010;
    16'b0000000000000000: out_v[323] = 10'b1000001100;
    16'b0000000000000001: out_v[323] = 10'b0110101000;
    16'b0010000000000010: out_v[323] = 10'b0001011101;
    16'b0001000000000011: out_v[323] = 10'b0111010001;
    16'b0011000000000110: out_v[323] = 10'b1000011111;
    16'b0000000000000110: out_v[323] = 10'b0110000101;
    16'b0010000000100001: out_v[323] = 10'b0000010110;
    16'b0011000000100000: out_v[323] = 10'b1101101110;
    16'b0001000000000001: out_v[323] = 10'b0110111000;
    16'b0001000000000101: out_v[323] = 10'b1101111010;
    16'b0011000000100010: out_v[323] = 10'b1010001111;
    16'b0001000000001100: out_v[323] = 10'b1110011011;
    16'b0010000000100000: out_v[323] = 10'b1001011010;
    16'b0010000000100010: out_v[323] = 10'b1110110110;
    16'b0101000000000000: out_v[323] = 10'b0000110001;
    16'b0011000000000101: out_v[323] = 10'b1001011110;
    16'b0001000100000000: out_v[323] = 10'b0011111011;
    16'b0001000100000001: out_v[323] = 10'b0001111111;
    16'b0011000000000100: out_v[323] = 10'b1011001000;
    16'b0000000000100000: out_v[323] = 10'b0101001010;
    16'b1001000000000000: out_v[323] = 10'b1100111001;
    16'b0011000000001100: out_v[323] = 10'b0101011010;
    16'b0011000100000010: out_v[323] = 10'b1110010100;
    16'b0100000000000011: out_v[323] = 10'b1010111000;
    16'b0100000000000010: out_v[323] = 10'b0110100011;
    16'b0111000100000010: out_v[323] = 10'b1010001010;
    16'b0110000000100010: out_v[323] = 10'b1101100111;
    16'b0011000100000110: out_v[323] = 10'b0010001001;
    16'b0011000100000011: out_v[323] = 10'b1000011110;
    16'b0011000001000011: out_v[323] = 10'b0101010111;
    16'b0110000000100011: out_v[323] = 10'b1101011101;
    16'b0100000000000000: out_v[323] = 10'b1010010001;
    16'b0111000000000100: out_v[323] = 10'b1111101100;
    16'b0101000000000100: out_v[323] = 10'b1111000111;
    16'b1101000000000000: out_v[323] = 10'b0011010110;
    16'b1100000000000000: out_v[323] = 10'b0000111010;
    16'b1111000000000000: out_v[323] = 10'b0111001111;
    16'b0111000001000011: out_v[323] = 10'b0010111010;
    16'b0111000010000011: out_v[323] = 10'b1010001111;
    16'b0110000000000110: out_v[323] = 10'b0010011011;
    16'b0010000000000111: out_v[323] = 10'b1110100011;
    16'b0111000000000110: out_v[323] = 10'b1111001011;
    16'b0110000000001001: out_v[323] = 10'b1011110010;
    16'b0110000000001101: out_v[323] = 10'b0101011111;
    16'b0111000000000101: out_v[323] = 10'b0001111011;
    16'b0010000000001101: out_v[323] = 10'b1100110110;
    16'b0110000000100000: out_v[323] = 10'b0111100110;
    16'b0010000000000101: out_v[323] = 10'b1111000000;
    16'b0111000000001101: out_v[323] = 10'b0111000110;
    16'b0110000000000101: out_v[323] = 10'b0011010110;
    16'b0000000000001101: out_v[323] = 10'b1101011010;
    16'b0010000000001001: out_v[323] = 10'b1001110110;
    16'b0011000000001101: out_v[323] = 10'b0010101111;
    16'b0001000001000011: out_v[323] = 10'b1000111001;
    16'b0100000001000011: out_v[323] = 10'b0111011111;
    16'b0000000001000011: out_v[323] = 10'b1011100010;
    16'b0101000001000011: out_v[323] = 10'b1010001010;
    16'b0001000001000010: out_v[323] = 10'b0011110011;
    16'b1000000000000001: out_v[323] = 10'b1000110111;
    16'b1001000000000001: out_v[323] = 10'b1101001110;
    default: out_v[323] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100010110000000: out_v[324] = 10'b1101110010;
    16'b0100010100000000: out_v[324] = 10'b0011100011;
    16'b0100110110000000: out_v[324] = 10'b1001110111;
    16'b0000010110000000: out_v[324] = 10'b0010011001;
    16'b0100000100000000: out_v[324] = 10'b0101110010;
    16'b0100100110000000: out_v[324] = 10'b0010100111;
    16'b0000000100000100: out_v[324] = 10'b0101100000;
    16'b0000000100000000: out_v[324] = 10'b0000110011;
    16'b0100010100000100: out_v[324] = 10'b1011100101;
    16'b0000010100000000: out_v[324] = 10'b1100111111;
    16'b0100010100000110: out_v[324] = 10'b0100010111;
    16'b0100010111000000: out_v[324] = 10'b0100110111;
    16'b0100000110000000: out_v[324] = 10'b0011011101;
    16'b0000100110000000: out_v[324] = 10'b0010011011;
    16'b0000000110000000: out_v[324] = 10'b1100010111;
    16'b0000110111000000: out_v[324] = 10'b0111111111;
    16'b0100000000000000: out_v[324] = 10'b0100101011;
    16'b0100000100000100: out_v[324] = 10'b1110111001;
    16'b0000010000000000: out_v[324] = 10'b1000000011;
    16'b0100000000000110: out_v[324] = 10'b0010110111;
    16'b0000000000000000: out_v[324] = 10'b1000000111;
    16'b0000110110000000: out_v[324] = 10'b0010010111;
    16'b0100010110000100: out_v[324] = 10'b0000111110;
    16'b0100010000000000: out_v[324] = 10'b0001001101;
    16'b0000000000000100: out_v[324] = 10'b0001010101;
    16'b0100000000000100: out_v[324] = 10'b0100100100;
    16'b0000010111000000: out_v[324] = 10'b0101010011;
    16'b0000000110000100: out_v[324] = 10'b0101011000;
    16'b0100010010000000: out_v[324] = 10'b0101100101;
    16'b0000010010000000: out_v[324] = 10'b0010011101;
    16'b0100010110000110: out_v[324] = 10'b1101001001;
    16'b0100000100000110: out_v[324] = 10'b1110010101;
    16'b0100000000000010: out_v[324] = 10'b1110101010;
    16'b0000000000000010: out_v[324] = 10'b0001110010;
    16'b0000000100000110: out_v[324] = 10'b0001110010;
    16'b0000000000000110: out_v[324] = 10'b0000111100;
    16'b0000010000000010: out_v[324] = 10'b0001011110;
    16'b0100010000000110: out_v[324] = 10'b0010110011;
    16'b0000000110000110: out_v[324] = 10'b1011000111;
    16'b0000010100000010: out_v[324] = 10'b1001110000;
    16'b0000010000000110: out_v[324] = 10'b0011001111;
    16'b0100010000000010: out_v[324] = 10'b0110100100;
    16'b0000010100000110: out_v[324] = 10'b0100110110;
    16'b0000000100000010: out_v[324] = 10'b1100100000;
    16'b0000000001000010: out_v[324] = 10'b1100011001;
    16'b0100000001000110: out_v[324] = 10'b1011000010;
    16'b0100000110000010: out_v[324] = 10'b1001001110;
    16'b0100000110000110: out_v[324] = 10'b1000100100;
    16'b0100000001000010: out_v[324] = 10'b1101011000;
    16'b0100000001000000: out_v[324] = 10'b0011111010;
    16'b0100010001000110: out_v[324] = 10'b1111011100;
    16'b0100000001000100: out_v[324] = 10'b1100011111;
    16'b0100010111000110: out_v[324] = 10'b1101110110;
    16'b0100000011000110: out_v[324] = 10'b0010110000;
    16'b0100000110000100: out_v[324] = 10'b1001001110;
    16'b0100000100000010: out_v[324] = 10'b1101011000;
    16'b0000000010000110: out_v[324] = 10'b1000110010;
    16'b0100000010000110: out_v[324] = 10'b0011111011;
    16'b0100000110100110: out_v[324] = 10'b1010101110;
    16'b0100000111000110: out_v[324] = 10'b1001111011;
    16'b0100010001000010: out_v[324] = 10'b0111011111;
    16'b0000000001000000: out_v[324] = 10'b1111100100;
    16'b0100000001100110: out_v[324] = 10'b1011001111;
    16'b0100000111100110: out_v[324] = 10'b0111010100;
    16'b0000000001000110: out_v[324] = 10'b1010000000;
    16'b0000000110000010: out_v[324] = 10'b0011101000;
    16'b0101000001000110: out_v[324] = 10'b1111111000;
    16'b0000000001000100: out_v[324] = 10'b0111001001;
    16'b0100010110000010: out_v[324] = 10'b1100001010;
    16'b0100000010000010: out_v[324] = 10'b0100011010;
    16'b0000010001000110: out_v[324] = 10'b0001100101;
    16'b0000010001000010: out_v[324] = 10'b1011011001;
    16'b0000010111000110: out_v[324] = 10'b0111110000;
    16'b0100010010000010: out_v[324] = 10'b1101010111;
    16'b0000010110000110: out_v[324] = 10'b1011111010;
    16'b0000010111000010: out_v[324] = 10'b0001010101;
    16'b0000010011000010: out_v[324] = 10'b0011110111;
    16'b1100010110000010: out_v[324] = 10'b0111010110;
    16'b0100010011000010: out_v[324] = 10'b0111110110;
    16'b0100010111000010: out_v[324] = 10'b1101100110;
    16'b0000010010000010: out_v[324] = 10'b0111000000;
    16'b0000010110000010: out_v[324] = 10'b0010011100;
    16'b0000010010000110: out_v[324] = 10'b0111000100;
    16'b0100010100000010: out_v[324] = 10'b0111011001;
    16'b1100010110000110: out_v[324] = 10'b1000110011;
    16'b0000010001000100: out_v[324] = 10'b1010011100;
    16'b0100010011000110: out_v[324] = 10'b1100110101;
    16'b0001010001000010: out_v[324] = 10'b0110101010;
    16'b0100010010000110: out_v[324] = 10'b0100000111;
    16'b0000010101000010: out_v[324] = 10'b0011001011;
    16'b0000010011000110: out_v[324] = 10'b1111110001;
    16'b0000010001000000: out_v[324] = 10'b0011110111;
    16'b0100010001000000: out_v[324] = 10'b1011001110;
    16'b1100010100000110: out_v[324] = 10'b0111110011;
    16'b0100100010000110: out_v[324] = 10'b1110001001;
    16'b0100100110000110: out_v[324] = 10'b1001000111;
    16'b0100000010000100: out_v[324] = 10'b0011010011;
    16'b0100100000000110: out_v[324] = 10'b0111110001;
    16'b0100100000000100: out_v[324] = 10'b0110010101;
    16'b0000010100000100: out_v[324] = 10'b0010110100;
    16'b0000010110000100: out_v[324] = 10'b1101101100;
    16'b0100010011000000: out_v[324] = 10'b0010100010;
    16'b1000010110000110: out_v[324] = 10'b1101011011;
    16'b0000110110000010: out_v[324] = 10'b1100110110;
    16'b1000010110000100: out_v[324] = 10'b0110101111;
    16'b0000000011000110: out_v[324] = 10'b0110010011;
    16'b0100000011000010: out_v[324] = 10'b1011010001;
    16'b0000000011000010: out_v[324] = 10'b0001100010;
    16'b0000000010000010: out_v[324] = 10'b0101100101;
    16'b0100000010000000: out_v[324] = 10'b1001000101;
    16'b0100000011000000: out_v[324] = 10'b1011101010;
    16'b1100110110000110: out_v[324] = 10'b0010110010;
    16'b1100000110000110: out_v[324] = 10'b0100001011;
    16'b1100010000000110: out_v[324] = 10'b1011000100;
    16'b1100010110000100: out_v[324] = 10'b0011011011;
    16'b1100000100000110: out_v[324] = 10'b0011111101;
    16'b0100100000000000: out_v[324] = 10'b0010000001;
    16'b1100000110000010: out_v[324] = 10'b0111101001;
    16'b0100110110000110: out_v[324] = 10'b0110011101;
    16'b0100100110000100: out_v[324] = 10'b0111010111;
    16'b1000010100000110: out_v[324] = 10'b1000001101;
    16'b0100100110000010: out_v[324] = 10'b1001011110;
    16'b1100000000000110: out_v[324] = 10'b1001000100;
    default: out_v[324] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000010101001: out_v[325] = 10'b0011011010;
    16'b0010000100101000: out_v[325] = 10'b1101001011;
    16'b0010000110101000: out_v[325] = 10'b1111010010;
    16'b0000000010001000: out_v[325] = 10'b1011100100;
    16'b0000100110100000: out_v[325] = 10'b1000011011;
    16'b0000100110101000: out_v[325] = 10'b1110011111;
    16'b0010000000101000: out_v[325] = 10'b1101001011;
    16'b0010000110101001: out_v[325] = 10'b1001100111;
    16'b1010000110101000: out_v[325] = 10'b1110101011;
    16'b0000000110001000: out_v[325] = 10'b0011001101;
    16'b0010100010101000: out_v[325] = 10'b0011101101;
    16'b0010000000001000: out_v[325] = 10'b0001100001;
    16'b0000000010101000: out_v[325] = 10'b0001110100;
    16'b0010000010001000: out_v[325] = 10'b1010100011;
    16'b0000000110101001: out_v[325] = 10'b0000110001;
    16'b1010000110100000: out_v[325] = 10'b1110111000;
    16'b0010000110001000: out_v[325] = 10'b1011001011;
    16'b0010000010100000: out_v[325] = 10'b1010110111;
    16'b0000000110101000: out_v[325] = 10'b1001100010;
    16'b0010000010101000: out_v[325] = 10'b1110010100;
    16'b0010100110101000: out_v[325] = 10'b1011000000;
    16'b0000000010001010: out_v[325] = 10'b1011110010;
    16'b0000100010000010: out_v[325] = 10'b0101011011;
    16'b0010000100001000: out_v[325] = 10'b1100110111;
    16'b0000000110001001: out_v[325] = 10'b0100101001;
    16'b0010000110001001: out_v[325] = 10'b0001010111;
    16'b0010000000100000: out_v[325] = 10'b1111110001;
    16'b0010000000000000: out_v[325] = 10'b1011100100;
    16'b0000000110001010: out_v[325] = 10'b0101101110;
    16'b0010100000000010: out_v[325] = 10'b1110001001;
    16'b0000000110000001: out_v[325] = 10'b0101000101;
    16'b0010100110101010: out_v[325] = 10'b1000111111;
    16'b0011000110000001: out_v[325] = 10'b1111100010;
    16'b0001000110000001: out_v[325] = 10'b0100110110;
    16'b0001000100000000: out_v[325] = 10'b0111001011;
    16'b0001000000000000: out_v[325] = 10'b1010000011;
    16'b0001000110000000: out_v[325] = 10'b1010111000;
    16'b0011000010000001: out_v[325] = 10'b1110010001;
    16'b0001000010000000: out_v[325] = 10'b1100010100;
    16'b0001000100000001: out_v[325] = 10'b0110001011;
    16'b0001000110000011: out_v[325] = 10'b1011010101;
    16'b0011000110100011: out_v[325] = 10'b1011100101;
    16'b0000000110100001: out_v[325] = 10'b1110000100;
    16'b0011000110000011: out_v[325] = 10'b0011110100;
    16'b0011000110100001: out_v[325] = 10'b1111100101;
    16'b0000000110000000: out_v[325] = 10'b0100111100;
    16'b0010000010000000: out_v[325] = 10'b0110100100;
    16'b0001000110100011: out_v[325] = 10'b1000111100;
    16'b0001000110100001: out_v[325] = 10'b1100110100;
    16'b0011000010100001: out_v[325] = 10'b1010011001;
    16'b0010000010000001: out_v[325] = 10'b1100101110;
    16'b0010000110100011: out_v[325] = 10'b1010101011;
    16'b0010000010100011: out_v[325] = 10'b1001101000;
    16'b0000000010100011: out_v[325] = 10'b1000011111;
    16'b0001000010100001: out_v[325] = 10'b1110010001;
    16'b0000000010100001: out_v[325] = 10'b1111010011;
    16'b0011000010000011: out_v[325] = 10'b1000010111;
    16'b0000000110000011: out_v[325] = 10'b0100100101;
    16'b0001000010000001: out_v[325] = 10'b0110000100;
    16'b0011000010100011: out_v[325] = 10'b0011100011;
    16'b0010000110100001: out_v[325] = 10'b1000011110;
    16'b0010000110000001: out_v[325] = 10'b0011100101;
    16'b0001000000000001: out_v[325] = 10'b0111000101;
    16'b0001000010000011: out_v[325] = 10'b1010110110;
    16'b0000000110100011: out_v[325] = 10'b1011100100;
    16'b0010000110000011: out_v[325] = 10'b1101110100;
    16'b0000000010000001: out_v[325] = 10'b0011000110;
    16'b0011000010100000: out_v[325] = 10'b0000111011;
    16'b0010000010000011: out_v[325] = 10'b1110110100;
    16'b0011000010000000: out_v[325] = 10'b1000111001;
    16'b0010000010100001: out_v[325] = 10'b0000011010;
    16'b0001000010100011: out_v[325] = 10'b0100000101;
    16'b0010000110000000: out_v[325] = 10'b1000011100;
    16'b0001000100100001: out_v[325] = 10'b0000101101;
    16'b0001100110000001: out_v[325] = 10'b1000100111;
    16'b0010000110100000: out_v[325] = 10'b0011010011;
    16'b0011000100101000: out_v[325] = 10'b1011010111;
    16'b0010000100000000: out_v[325] = 10'b1101100001;
    16'b0000000100100000: out_v[325] = 10'b0101011010;
    16'b0010000100001010: out_v[325] = 10'b0000111100;
    16'b0000000100101000: out_v[325] = 10'b1011000110;
    16'b0010000100100000: out_v[325] = 10'b1111001010;
    16'b0001000100100000: out_v[325] = 10'b1101001101;
    16'b0011000000000000: out_v[325] = 10'b0000100111;
    16'b0011000100000000: out_v[325] = 10'b1011110111;
    16'b0011000110100000: out_v[325] = 10'b0101011011;
    16'b0011000100100001: out_v[325] = 10'b0001011001;
    16'b0001000100101000: out_v[325] = 10'b0100011001;
    16'b0011000110000000: out_v[325] = 10'b0000111000;
    16'b0011000100001010: out_v[325] = 10'b1101011011;
    16'b0010000100000010: out_v[325] = 10'b0110011111;
    16'b0010000110001010: out_v[325] = 10'b0011011101;
    16'b0000000110100000: out_v[325] = 10'b1000011010;
    16'b0011000100100000: out_v[325] = 10'b1001010010;
    16'b0011000000101000: out_v[325] = 10'b0011001010;
    16'b0000000110000010: out_v[325] = 10'b1001011011;
    16'b0000000100000000: out_v[325] = 10'b1101010100;
    16'b0000000000100000: out_v[325] = 10'b0011110110;
    16'b0011000000100000: out_v[325] = 10'b0100011011;
    16'b0011000000100001: out_v[325] = 10'b1100010011;
    16'b0011000110101000: out_v[325] = 10'b1011101001;
    16'b0001000110101000: out_v[325] = 10'b0101000001;
    16'b0001000110100000: out_v[325] = 10'b0000011011;
    16'b0001000000101001: out_v[325] = 10'b0010111011;
    16'b0000000100101001: out_v[325] = 10'b1000111110;
    16'b0001000000001100: out_v[325] = 10'b1000011011;
    16'b0001000010001001: out_v[325] = 10'b0110100011;
    16'b0001000110001000: out_v[325] = 10'b1001110010;
    16'b0001000000001000: out_v[325] = 10'b1000010001;
    16'b0011000010001000: out_v[325] = 10'b1001011110;
    16'b0001000010001000: out_v[325] = 10'b0101110111;
    16'b0001000100001001: out_v[325] = 10'b1000010101;
    16'b0001000110001001: out_v[325] = 10'b0111000101;
    16'b0001000000001001: out_v[325] = 10'b0010101101;
    16'b0000000000001000: out_v[325] = 10'b1101010100;
    16'b0001000100001000: out_v[325] = 10'b0001010111;
    16'b0011000010001001: out_v[325] = 10'b0100011000;
    16'b0000000000101000: out_v[325] = 10'b1100110001;
    16'b0000000100001001: out_v[325] = 10'b1000111001;
    16'b0000000000101001: out_v[325] = 10'b1000111000;
    16'b0000000000100001: out_v[325] = 10'b0010111001;
    16'b0000000010001001: out_v[325] = 10'b1011001110;
    16'b0001000100101001: out_v[325] = 10'b0010111010;
    16'b0001000000101000: out_v[325] = 10'b1000100001;
    16'b0000000100001000: out_v[325] = 10'b1011000010;
    16'b0000000000001001: out_v[325] = 10'b0100111110;
    16'b0001000000100001: out_v[325] = 10'b0011101101;
    16'b0001000100101011: out_v[325] = 10'b1100001101;
    16'b0001000000001101: out_v[325] = 10'b0011101111;
    16'b0000000000000001: out_v[325] = 10'b1000011110;
    16'b0000000100000001: out_v[325] = 10'b1010110000;
    16'b0011000110001000: out_v[325] = 10'b1000101000;
    16'b0000000010000000: out_v[325] = 10'b1101101010;
    16'b0010000000001010: out_v[325] = 10'b1111110000;
    16'b0010000100001001: out_v[325] = 10'b1001111011;
    16'b0010000010001010: out_v[325] = 10'b1010100100;
    16'b0011000100001000: out_v[325] = 10'b0011100111;
    16'b0001000010101000: out_v[325] = 10'b0010101111;
    16'b0000000000000000: out_v[325] = 10'b1011011100;
    16'b0011000000001000: out_v[325] = 10'b1111000100;
    16'b0000000000001010: out_v[325] = 10'b0001001100;
    16'b0000000100001101: out_v[325] = 10'b1001100111;
    16'b0000000010100000: out_v[325] = 10'b0000110101;
    16'b0011000010101000: out_v[325] = 10'b1001000100;
    16'b0001000010101011: out_v[325] = 10'b1111010011;
    16'b0001000010101001: out_v[325] = 10'b0111001111;
    16'b0001100010101001: out_v[325] = 10'b1111110001;
    16'b0001000110101001: out_v[325] = 10'b0111101100;
    16'b0000100010101000: out_v[325] = 10'b1001011100;
    16'b0001000010001011: out_v[325] = 10'b1001001010;
    16'b0011000010101001: out_v[325] = 10'b1110001000;
    16'b0000100010101001: out_v[325] = 10'b1111100010;
    16'b0011000110101001: out_v[325] = 10'b1101011010;
    16'b0000000010001011: out_v[325] = 10'b0011100011;
    16'b0000000000000100: out_v[325] = 10'b0000001111;
    16'b0000000100000100: out_v[325] = 10'b0100110101;
    16'b0000000110000100: out_v[325] = 10'b0110111011;
    16'b0000000100001100: out_v[325] = 10'b0111001100;
    16'b0000001100000000: out_v[325] = 10'b1101111011;
    16'b0001000100000100: out_v[325] = 10'b1001111100;
    16'b0001000110000100: out_v[325] = 10'b1011110001;
    16'b0000001100000100: out_v[325] = 10'b0011010111;
    16'b0000000100101100: out_v[325] = 10'b0111001111;
    16'b0001000100001100: out_v[325] = 10'b0001110011;
    16'b0000000110001100: out_v[325] = 10'b0011001010;
    16'b0000001100100000: out_v[325] = 10'b1000110110;
    16'b0001000110000101: out_v[325] = 10'b0111010011;
    16'b0001000100000101: out_v[325] = 10'b0011101001;
    16'b0000000100100100: out_v[325] = 10'b0101011011;
    16'b0001000110001100: out_v[325] = 10'b0010001001;
    16'b0011000110001001: out_v[325] = 10'b1110000100;
    16'b0011000000000001: out_v[325] = 10'b0001111010;
    16'b0011000000001001: out_v[325] = 10'b0011010111;
    16'b0011000100000001: out_v[325] = 10'b0101000001;
    16'b0001000110101011: out_v[325] = 10'b0100100110;
    16'b0011000100001001: out_v[325] = 10'b0110110111;
    16'b0001000110001011: out_v[325] = 10'b0110010011;
    16'b0010000000000001: out_v[325] = 10'b0100000110;
    16'b0011000000101001: out_v[325] = 10'b0110100000;
    16'b0000000000001100: out_v[325] = 10'b0010111110;
    16'b0001000010001100: out_v[325] = 10'b0000011111;
    16'b0001000100001101: out_v[325] = 10'b1001000110;
    16'b0001000110001101: out_v[325] = 10'b1101000110;
    16'b0000000100100001: out_v[325] = 10'b1011101010;
    default: out_v[325] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000001001000010: out_v[326] = 10'b0100101000;
    16'b0000010001001010: out_v[326] = 10'b1101000100;
    16'b0000011001001010: out_v[326] = 10'b0000100101;
    16'b0000000001000010: out_v[326] = 10'b0100110111;
    16'b0000000001001010: out_v[326] = 10'b1001101101;
    16'b0000000001001000: out_v[326] = 10'b1110010111;
    16'b1000001001001010: out_v[326] = 10'b0011100110;
    16'b0000011000001010: out_v[326] = 10'b0111101010;
    16'b1000001001000010: out_v[326] = 10'b1000101100;
    16'b0000001001001010: out_v[326] = 10'b0111000010;
    16'b0000001000000000: out_v[326] = 10'b1100100011;
    16'b0000001001000000: out_v[326] = 10'b1111011000;
    16'b0000010000000010: out_v[326] = 10'b0110100001;
    16'b0000001000001010: out_v[326] = 10'b0100011111;
    16'b0000010000001010: out_v[326] = 10'b0111011001;
    16'b0000001001001000: out_v[326] = 10'b1010011110;
    16'b0000001000000010: out_v[326] = 10'b0001100011;
    16'b0000001000001000: out_v[326] = 10'b0011111001;
    16'b0000011000001000: out_v[326] = 10'b1101010001;
    16'b1000000001000010: out_v[326] = 10'b0111100001;
    16'b1000011001001010: out_v[326] = 10'b0001110111;
    16'b0000010001000010: out_v[326] = 10'b1100110110;
    16'b0000000000001000: out_v[326] = 10'b1010110000;
    16'b0000000000001010: out_v[326] = 10'b0110110001;
    16'b1000000001001010: out_v[326] = 10'b1111011001;
    16'b0000011000000010: out_v[326] = 10'b1011110100;
    16'b0000011001000010: out_v[326] = 10'b1000111110;
    16'b0000000001000000: out_v[326] = 10'b0010010110;
    16'b0000000000000010: out_v[326] = 10'b0100111010;
    16'b0000010000001000: out_v[326] = 10'b1100000001;
    16'b1000001000001010: out_v[326] = 10'b1111000001;
    16'b1000000000000010: out_v[326] = 10'b1111010011;
    16'b0000000000000000: out_v[326] = 10'b1011000010;
    16'b0000010001000000: out_v[326] = 10'b0011001110;
    16'b1000000000000000: out_v[326] = 10'b0101110010;
    16'b0000010000000000: out_v[326] = 10'b0110111000;
    16'b0000011001000000: out_v[326] = 10'b0111011000;
    16'b1000001001000000: out_v[326] = 10'b1011001111;
    16'b1000011001000010: out_v[326] = 10'b0100110110;
    16'b0000011000000000: out_v[326] = 10'b1010011100;
    16'b1000011000000010: out_v[326] = 10'b1011100111;
    16'b1000001000000000: out_v[326] = 10'b0110000101;
    16'b1000001000000010: out_v[326] = 10'b0011001110;
    16'b0000100001000000: out_v[326] = 10'b0100011011;
    16'b0000110001000000: out_v[326] = 10'b1001100111;
    16'b0000110000000000: out_v[326] = 10'b0001111110;
    16'b0000010001001000: out_v[326] = 10'b1010110100;
    16'b1000000001000000: out_v[326] = 10'b1111011011;
    16'b0000100000000010: out_v[326] = 10'b1011010101;
    16'b0000100000001010: out_v[326] = 10'b1010101000;
    16'b1000000001001000: out_v[326] = 10'b1010010000;
    16'b1000000000001010: out_v[326] = 10'b1101010011;
    16'b1000000000001000: out_v[326] = 10'b1011110000;
    16'b1000010001001000: out_v[326] = 10'b1011111100;
    16'b0000000000010010: out_v[326] = 10'b1110001101;
    16'b0000000001010010: out_v[326] = 10'b1010111111;
    16'b0000000000011010: out_v[326] = 10'b0000110110;
    16'b0000000001011010: out_v[326] = 10'b0000101000;
    16'b0000000000010000: out_v[326] = 10'b0001111001;
    16'b0000100000000000: out_v[326] = 10'b0111111010;
    16'b1000011000001010: out_v[326] = 10'b1100110010;
    16'b0000100001001010: out_v[326] = 10'b1111001010;
    16'b0000000001001001: out_v[326] = 10'b0110110111;
    16'b0000100001000010: out_v[326] = 10'b1111000011;
    16'b0000000001000001: out_v[326] = 10'b1011000011;
    16'b0000110000000010: out_v[326] = 10'b1010110111;
    16'b0000110001000010: out_v[326] = 10'b0110101001;
    16'b0000100001001000: out_v[326] = 10'b1111110110;
    default: out_v[326] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010001000000101: out_v[327] = 10'b0011001011;
    16'b0011000001000100: out_v[327] = 10'b0111100000;
    16'b0010000000000101: out_v[327] = 10'b0010110110;
    16'b0011000000000101: out_v[327] = 10'b1100110000;
    16'b0010001000000100: out_v[327] = 10'b0001010010;
    16'b0010010000000101: out_v[327] = 10'b1100110101;
    16'b0010000001000100: out_v[327] = 10'b1110011111;
    16'b0010000001000101: out_v[327] = 10'b0000011110;
    16'b0000000000000101: out_v[327] = 10'b1010100001;
    16'b0010011000000100: out_v[327] = 10'b0001011110;
    16'b0000011000000101: out_v[327] = 10'b1101010110;
    16'b0010000000000100: out_v[327] = 10'b0001000101;
    16'b0010001000000000: out_v[327] = 10'b1101010101;
    16'b0010011000000101: out_v[327] = 10'b0001010101;
    16'b0000000000000000: out_v[327] = 10'b0010000011;
    16'b0000000000000001: out_v[327] = 10'b0000100010;
    16'b0000001000000101: out_v[327] = 10'b0110011000;
    16'b0010010000000100: out_v[327] = 10'b1011010010;
    16'b0010001001000101: out_v[327] = 10'b1010100011;
    16'b0011000001000101: out_v[327] = 10'b1001110001;
    16'b0000001000000000: out_v[327] = 10'b0101000101;
    16'b0011010001000100: out_v[327] = 10'b1010011101;
    16'b0010001001000100: out_v[327] = 10'b1110000101;
    16'b0000001000000001: out_v[327] = 10'b0101001000;
    16'b0000000001000001: out_v[327] = 10'b1001000111;
    16'b0010010001000101: out_v[327] = 10'b1000101110;
    16'b0000000001000000: out_v[327] = 10'b0000111011;
    16'b0000000001000101: out_v[327] = 10'b0111000000;
    16'b0000010000000101: out_v[327] = 10'b1110101011;
    16'b0000000000000100: out_v[327] = 10'b1001000111;
    16'b0011000000000100: out_v[327] = 10'b1101001111;
    16'b0000001000000100: out_v[327] = 10'b0001110011;
    16'b0000011001000000: out_v[327] = 10'b0010011011;
    16'b0000011000000000: out_v[327] = 10'b0100110111;
    16'b0000010000000000: out_v[327] = 10'b0000111010;
    16'b0001011000000000: out_v[327] = 10'b0111010010;
    16'b0001011001000000: out_v[327] = 10'b0100110111;
    16'b0000010000000001: out_v[327] = 10'b1011110100;
    16'b0000011000000100: out_v[327] = 10'b0100001010;
    16'b0011001001000101: out_v[327] = 10'b0001011110;
    16'b0000001001000000: out_v[327] = 10'b1001010101;
    16'b0011001000000101: out_v[327] = 10'b0000000110;
    16'b0010000000000000: out_v[327] = 10'b1110101101;
    16'b0011001000000100: out_v[327] = 10'b0111100011;
    16'b0011011000000101: out_v[327] = 10'b1111100100;
    16'b0001001000000000: out_v[327] = 10'b0011011010;
    16'b0000011000000001: out_v[327] = 10'b1110010100;
    16'b0010011001000100: out_v[327] = 10'b1001001011;
    16'b0010011000000000: out_v[327] = 10'b1110110100;
    16'b0011011000000100: out_v[327] = 10'b1110111111;
    16'b0001001001000001: out_v[327] = 10'b0100010100;
    16'b0001001001000000: out_v[327] = 10'b1111000000;
    16'b0011010000000101: out_v[327] = 10'b0011011010;
    16'b0001010000000100: out_v[327] = 10'b1110111011;
    16'b0000010000000100: out_v[327] = 10'b1011011010;
    16'b0011010000000100: out_v[327] = 10'b0111100001;
    16'b0010010000000001: out_v[327] = 10'b1111011011;
    16'b0010010000000000: out_v[327] = 10'b1101011011;
    16'b0011010001000000: out_v[327] = 10'b1100101011;
    16'b0001010000000000: out_v[327] = 10'b0001001100;
    16'b0011010000000000: out_v[327] = 10'b0111111110;
    16'b0010010001000100: out_v[327] = 10'b0100011010;
    16'b0011010001000101: out_v[327] = 10'b0111001110;
    16'b0001010001000000: out_v[327] = 10'b0001111010;
    16'b0001010000000101: out_v[327] = 10'b1010011110;
    16'b0010011000000001: out_v[327] = 10'b1000111101;
    16'b0000010001000001: out_v[327] = 10'b1110001011;
    16'b0100000000000001: out_v[327] = 10'b1011110011;
    16'b0010000000000001: out_v[327] = 10'b1000100010;
    16'b0100000000000000: out_v[327] = 10'b0011111011;
    16'b0000010001000000: out_v[327] = 10'b1100010100;
    16'b0000011001000001: out_v[327] = 10'b0110010100;
    16'b0000001001000001: out_v[327] = 10'b0011010100;
    16'b0010000001000001: out_v[327] = 10'b1011001011;
    16'b0010001000000001: out_v[327] = 10'b1111001111;
    16'b0110000001000101: out_v[327] = 10'b1100110000;
    16'b0000010001000101: out_v[327] = 10'b1110011010;
    16'b0001000001000000: out_v[327] = 10'b1010101001;
    16'b0100000001000000: out_v[327] = 10'b0110100011;
    16'b0100000001000001: out_v[327] = 10'b0011101110;
    16'b0010000001000000: out_v[327] = 10'b1011000101;
    16'b0010010010000101: out_v[327] = 10'b1010110010;
    16'b0001011000000001: out_v[327] = 10'b1011110101;
    16'b0001000000000001: out_v[327] = 10'b1110000001;
    16'b0001001000000001: out_v[327] = 10'b0101101010;
    16'b0010011001000101: out_v[327] = 10'b1101000011;
    16'b0010011001000001: out_v[327] = 10'b1100000100;
    16'b0001011001000001: out_v[327] = 10'b0010010100;
    default: out_v[327] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000010000000010: out_v[328] = 10'b0010010111;
    16'b1110010000000010: out_v[328] = 10'b0101100111;
    16'b1010000010000010: out_v[328] = 10'b0111111001;
    16'b0010010000000010: out_v[328] = 10'b1010001011;
    16'b1000010000000011: out_v[328] = 10'b1100110110;
    16'b1010000010000011: out_v[328] = 10'b1010010111;
    16'b1000000000000010: out_v[328] = 10'b1000100000;
    16'b1010010000000010: out_v[328] = 10'b0011001011;
    16'b1010000000000010: out_v[328] = 10'b1001011010;
    16'b1001010000000011: out_v[328] = 10'b1011111100;
    16'b1010000000100000: out_v[328] = 10'b1101110101;
    16'b1011010000000010: out_v[328] = 10'b0001111010;
    16'b0010010000000011: out_v[328] = 10'b1001110011;
    16'b1010010000000011: out_v[328] = 10'b1111001101;
    16'b1110010000000011: out_v[328] = 10'b0011111110;
    16'b1010010000100000: out_v[328] = 10'b1011000111;
    16'b1010001000100000: out_v[328] = 10'b1011011111;
    16'b1001010000000001: out_v[328] = 10'b1111000001;
    16'b0010010000100010: out_v[328] = 10'b0100001111;
    16'b1000000000100000: out_v[328] = 10'b1110001011;
    16'b1011010000000011: out_v[328] = 10'b0010000111;
    16'b1010010000100010: out_v[328] = 10'b1110010010;
    16'b1111010000000011: out_v[328] = 10'b0011011111;
    16'b1000001000100000: out_v[328] = 10'b1110100011;
    16'b1010000000000011: out_v[328] = 10'b1101000011;
    16'b0010010000100000: out_v[328] = 10'b0010001011;
    16'b1111010000000010: out_v[328] = 10'b0001110011;
    16'b1010000010100010: out_v[328] = 10'b1001111110;
    16'b1011000000000011: out_v[328] = 10'b0100101110;
    16'b1011000010000010: out_v[328] = 10'b1011001101;
    16'b1110000000000010: out_v[328] = 10'b1001010111;
    16'b1000010000000010: out_v[328] = 10'b0101001111;
    16'b1010000010100000: out_v[328] = 10'b0111011011;
    16'b1000000000000000: out_v[328] = 10'b0011100101;
    16'b1011000000000010: out_v[328] = 10'b1101111010;
    16'b0000010000000011: out_v[328] = 10'b1000010010;
    16'b1010011000100000: out_v[328] = 10'b1100110011;
    16'b1000010000000001: out_v[328] = 10'b0011000101;
    16'b1010000000100010: out_v[328] = 10'b1011011100;
    16'b1001000000000000: out_v[328] = 10'b0110110001;
    16'b0001000000000000: out_v[328] = 10'b1010110100;
    16'b0001000000000001: out_v[328] = 10'b1101001001;
    16'b1101000000000000: out_v[328] = 10'b0101110101;
    16'b0101000000000000: out_v[328] = 10'b1000111110;
    16'b1001000000000001: out_v[328] = 10'b1011101000;
    16'b1001010000000000: out_v[328] = 10'b0010010110;
    16'b0000000000000000: out_v[328] = 10'b0101001010;
    16'b0000000000000001: out_v[328] = 10'b0110010111;
    16'b1001000000100000: out_v[328] = 10'b1011011011;
    16'b0001001000100000: out_v[328] = 10'b0011110100;
    16'b1010010000000001: out_v[328] = 10'b0100011011;
    16'b1000000000000001: out_v[328] = 10'b1100110110;
    16'b1000010000100011: out_v[328] = 10'b0101001010;
    16'b1001010000100000: out_v[328] = 10'b1000100110;
    16'b1000000000100011: out_v[328] = 10'b1101110100;
    16'b0000000000000011: out_v[328] = 10'b0111100101;
    16'b1000011000100011: out_v[328] = 10'b1101101101;
    16'b1010010000100011: out_v[328] = 10'b0101000100;
    16'b1000000000100001: out_v[328] = 10'b0011010111;
    16'b1000001000000000: out_v[328] = 10'b1000100111;
    16'b1010011000000011: out_v[328] = 10'b1100010110;
    16'b1000010000100001: out_v[328] = 10'b1011101100;
    16'b1001011000100000: out_v[328] = 10'b0111110101;
    16'b1000011000000011: out_v[328] = 10'b1101110111;
    16'b0001011000000011: out_v[328] = 10'b0111110011;
    16'b0001010000000011: out_v[328] = 10'b1001111001;
    16'b1001001000100000: out_v[328] = 10'b0101001000;
    16'b1000001000100001: out_v[328] = 10'b1110011001;
    16'b1001000000100001: out_v[328] = 10'b1110110110;
    16'b1001011000100011: out_v[328] = 10'b0011001111;
    16'b1001010000100011: out_v[328] = 10'b1111010011;
    16'b1001010000100001: out_v[328] = 10'b0100010000;
    16'b1000001000000011: out_v[328] = 10'b1000110111;
    16'b0001000000100000: out_v[328] = 10'b1011001111;
    16'b1010011000100011: out_v[328] = 10'b0100100110;
    16'b0000010000000001: out_v[328] = 10'b1001100110;
    16'b0001000000000011: out_v[328] = 10'b1010010010;
    16'b0001010000000001: out_v[328] = 10'b1100100011;
    16'b1001000000000011: out_v[328] = 10'b0110100010;
    16'b0001010000100000: out_v[328] = 10'b1001111100;
    16'b1000000000000011: out_v[328] = 10'b1001111100;
    16'b1000010000000000: out_v[328] = 10'b0101010100;
    16'b0000010000100011: out_v[328] = 10'b0011101100;
    16'b0001010000100011: out_v[328] = 10'b1100000011;
    16'b1101001000000010: out_v[328] = 10'b1111011110;
    16'b1001000000000010: out_v[328] = 10'b0001001111;
    16'b1001001000000010: out_v[328] = 10'b1011101110;
    16'b1001001000000011: out_v[328] = 10'b0001111010;
    16'b0001000000000010: out_v[328] = 10'b0100000010;
    16'b0001010000000010: out_v[328] = 10'b0011001110;
    16'b0001001000000010: out_v[328] = 10'b0101000010;
    16'b0101000000000010: out_v[328] = 10'b0111001011;
    16'b1001010000000010: out_v[328] = 10'b0000100111;
    16'b1101000000000011: out_v[328] = 10'b1001110101;
    16'b0001001000000011: out_v[328] = 10'b0011011011;
    16'b0001001000100010: out_v[328] = 10'b1111010011;
    16'b1011001000100000: out_v[328] = 10'b1011000100;
    16'b1101001000000011: out_v[328] = 10'b0101110111;
    16'b0101000000000001: out_v[328] = 10'b1000101000;
    16'b1101000000000001: out_v[328] = 10'b1110100101;
    16'b0101001000000010: out_v[328] = 10'b1111110001;
    16'b1001001000100010: out_v[328] = 10'b0111111001;
    16'b0001001000100011: out_v[328] = 10'b0101011011;
    16'b1101000000000010: out_v[328] = 10'b0011110010;
    16'b1011001000000010: out_v[328] = 10'b0011011011;
    16'b1001000000100010: out_v[328] = 10'b0001110001;
    16'b0101000000000011: out_v[328] = 10'b0101110111;
    16'b1101010000000010: out_v[328] = 10'b1110100010;
    16'b0001001000000001: out_v[328] = 10'b1100010100;
    16'b0101010000000011: out_v[328] = 10'b0001101011;
    16'b1011001000100010: out_v[328] = 10'b1011100010;
    16'b0101010000000010: out_v[328] = 10'b0000011110;
    16'b0001010000000000: out_v[328] = 10'b1010101100;
    16'b0010000000000001: out_v[328] = 10'b1100011001;
    16'b0011010000000001: out_v[328] = 10'b0100111000;
    16'b0010011000100011: out_v[328] = 10'b0100011110;
    16'b0000011000000001: out_v[328] = 10'b0111001011;
    16'b0010010000000001: out_v[328] = 10'b0001101001;
    16'b0000010000000000: out_v[328] = 10'b1101110000;
    16'b0010011000000011: out_v[328] = 10'b0001100111;
    16'b0011010000000011: out_v[328] = 10'b1001000111;
    16'b0000011000000011: out_v[328] = 10'b1010100101;
    16'b0011000000000001: out_v[328] = 10'b0000011001;
    16'b0010010010000011: out_v[328] = 10'b1001101010;
    16'b0000010010000011: out_v[328] = 10'b0011010001;
    16'b1100000000000011: out_v[328] = 10'b1111010110;
    16'b0000000000000010: out_v[328] = 10'b1011110111;
    16'b0100000000000001: out_v[328] = 10'b1110010010;
    16'b1100000000000001: out_v[328] = 10'b1011010110;
    16'b1011000000100000: out_v[328] = 10'b0001111001;
    16'b1000000000100010: out_v[328] = 10'b1111100111;
    16'b1100010000000001: out_v[328] = 10'b0101001111;
    16'b0100000000000010: out_v[328] = 10'b0001110110;
    16'b0000000000100010: out_v[328] = 10'b0001001011;
    16'b0100010000000001: out_v[328] = 10'b1000001100;
    16'b0100000000000011: out_v[328] = 10'b0100011001;
    16'b0000010000100010: out_v[328] = 10'b0011110011;
    16'b0010010000000000: out_v[328] = 10'b0001100110;
    16'b0010010000100001: out_v[328] = 10'b1111100010;
    16'b0010000000000011: out_v[328] = 10'b1100011110;
    16'b0010010000100011: out_v[328] = 10'b0110111111;
    16'b0000010000100000: out_v[328] = 10'b0100110111;
    16'b0011010000000010: out_v[328] = 10'b1001101000;
    16'b0011010000100000: out_v[328] = 10'b1011000011;
    16'b0000001000000001: out_v[328] = 10'b0100101111;
    16'b0111000000000001: out_v[328] = 10'b0011101111;
    16'b0011000000000010: out_v[328] = 10'b0101110001;
    16'b0000000000001001: out_v[328] = 10'b0111100110;
    16'b0000001000000011: out_v[328] = 10'b1100011101;
    16'b0000001000001001: out_v[328] = 10'b0110111011;
    16'b0001000000001001: out_v[328] = 10'b0011001111;
    16'b0011000000000011: out_v[328] = 10'b0110001110;
    16'b1100000000000000: out_v[328] = 10'b1111010000;
    16'b0011001000000011: out_v[328] = 10'b1100110111;
    16'b0110000000000001: out_v[328] = 10'b1001111100;
    16'b0100000000000000: out_v[328] = 10'b0010111001;
    16'b0100001000000001: out_v[328] = 10'b1101100011;
    16'b1110000000000001: out_v[328] = 10'b0101011011;
    16'b1010010000000000: out_v[328] = 10'b0110001000;
    16'b1101010000000000: out_v[328] = 10'b0100100111;
    16'b1100010000000000: out_v[328] = 10'b1001010111;
    16'b1110010000000001: out_v[328] = 10'b1101001011;
    16'b1101010000000001: out_v[328] = 10'b1101000110;
    16'b1010000000000001: out_v[328] = 10'b0001001011;
    16'b1110010000000000: out_v[328] = 10'b0111011110;
    16'b0110010000000001: out_v[328] = 10'b1010100010;
    default: out_v[328] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000001110000: out_v[329] = 10'b0101110110;
    16'b0000101001111110: out_v[329] = 10'b0111011101;
    16'b0001100000111110: out_v[329] = 10'b1001111111;
    16'b0001100001111110: out_v[329] = 10'b0110111111;
    16'b0000000001111000: out_v[329] = 10'b1000110101;
    16'b0000000001111100: out_v[329] = 10'b0001011110;
    16'b0001101000111110: out_v[329] = 10'b1111001111;
    16'b0001101001111110: out_v[329] = 10'b0100000001;
    16'b0000000000111000: out_v[329] = 10'b1001001111;
    16'b0000100001111100: out_v[329] = 10'b0011001010;
    16'b0000000000111100: out_v[329] = 10'b0110100111;
    16'b0000000000101100: out_v[329] = 10'b1010011001;
    16'b0000000010111000: out_v[329] = 10'b1100110011;
    16'b0001100001111100: out_v[329] = 10'b1010110011;
    16'b0001101001110110: out_v[329] = 10'b1000111011;
    16'b0000100011111110: out_v[329] = 10'b0100010011;
    16'b0000100000111100: out_v[329] = 10'b0101010111;
    16'b0000000000011100: out_v[329] = 10'b0001110011;
    16'b0000100010111100: out_v[329] = 10'b1011011011;
    16'b0000100000111110: out_v[329] = 10'b0111001010;
    16'b0000100001111110: out_v[329] = 10'b0111111011;
    16'b0001100011111110: out_v[329] = 10'b0100010011;
    16'b0000000011111100: out_v[329] = 10'b0101010101;
    16'b0001101001110010: out_v[329] = 10'b0101001011;
    16'b0001101001011110: out_v[329] = 10'b0111000001;
    16'b0001100000111100: out_v[329] = 10'b0100110011;
    16'b0000000001111110: out_v[329] = 10'b1111001110;
    16'b0000000001010000: out_v[329] = 10'b0001000011;
    16'b0001101000011110: out_v[329] = 10'b1101000001;
    16'b0000001001111110: out_v[329] = 10'b0101001011;
    16'b0001100000110010: out_v[329] = 10'b0011011011;
    16'b0001100001110110: out_v[329] = 10'b1111011110;
    16'b0000101011111110: out_v[329] = 10'b1010010011;
    16'b0000101001111100: out_v[329] = 10'b0011001111;
    16'b0000000010111100: out_v[329] = 10'b1001010001;
    16'b0000101001011110: out_v[329] = 10'b1010111111;
    16'b0001101001111100: out_v[329] = 10'b0111000111;
    16'b0000000000100000: out_v[329] = 10'b1011101111;
    16'b0000100011111100: out_v[329] = 10'b1111110110;
    16'b0000000000110000: out_v[329] = 10'b1100000010;
    16'b0001100000110110: out_v[329] = 10'b0000111110;
    16'b0001101001101110: out_v[329] = 10'b1010100100;
    16'b0001101011111110: out_v[329] = 10'b1110110111;
    16'b0000000011111000: out_v[329] = 10'b1110111011;
    16'b0001100000101110: out_v[329] = 10'b0110111010;
    16'b0000100001011100: out_v[329] = 10'b0111000001;
    16'b0000001001010000: out_v[329] = 10'b1011100011;
    16'b0000000000000000: out_v[329] = 10'b0111001111;
    16'b0000000010000000: out_v[329] = 10'b1111101000;
    16'b0000000001000000: out_v[329] = 10'b1001010011;
    16'b0000001000010000: out_v[329] = 10'b0101000110;
    16'b0000000000010000: out_v[329] = 10'b0110001110;
    16'b0000001000000000: out_v[329] = 10'b0010100011;
    16'b0000000010100000: out_v[329] = 10'b0111000011;
    16'b0000000010010000: out_v[329] = 10'b1001001100;
    16'b0000100011011100: out_v[329] = 10'b0100110111;
    16'b0000000011010000: out_v[329] = 10'b1011011110;
    16'b0000000011000000: out_v[329] = 10'b1110110100;
    16'b0000100011010000: out_v[329] = 10'b0011110000;
    16'b0000100000101100: out_v[329] = 10'b0001010110;
    16'b0000100011110000: out_v[329] = 10'b0011100110;
    16'b0001101011011110: out_v[329] = 10'b0010111110;
    16'b0001101001001110: out_v[329] = 10'b0010001110;
    16'b0001100001001100: out_v[329] = 10'b0011010011;
    16'b0000100000000000: out_v[329] = 10'b0101011110;
    16'b0000000010110000: out_v[329] = 10'b1001100111;
    16'b0001100011011100: out_v[329] = 10'b1110010010;
    16'b0001100011001100: out_v[329] = 10'b1010000011;
    16'b0000100011001100: out_v[329] = 10'b0100100100;
    16'b0000100000001100: out_v[329] = 10'b1100110111;
    16'b0010000000010000: out_v[329] = 10'b1101100101;
    16'b0001100000001100: out_v[329] = 10'b1000100100;
    16'b0000100010010000: out_v[329] = 10'b0010010101;
    16'b0000000011110000: out_v[329] = 10'b0000100100;
    16'b0000101001110000: out_v[329] = 10'b1110011100;
    16'b0000100000100000: out_v[329] = 10'b0000110110;
    16'b0001100000101100: out_v[329] = 10'b0010100100;
    16'b0001101001001100: out_v[329] = 10'b1011010100;
    16'b0010000011010000: out_v[329] = 10'b0111110011;
    16'b0010000000000000: out_v[329] = 10'b0111110011;
    16'b0010000010010000: out_v[329] = 10'b1101110010;
    16'b0000100011000000: out_v[329] = 10'b0011110011;
    16'b0000100001110000: out_v[329] = 10'b1010011110;
    16'b0001100001101100: out_v[329] = 10'b0111110110;
    16'b0001100011000000: out_v[329] = 10'b0110100111;
    16'b0000000000001100: out_v[329] = 10'b1000111010;
    16'b0001101011001110: out_v[329] = 10'b1000101111;
    16'b0000100001010000: out_v[329] = 10'b1011011100;
    16'b0000000000001000: out_v[329] = 10'b1011100110;
    16'b0000000000011000: out_v[329] = 10'b1110110110;
    16'b0001100011010000: out_v[329] = 10'b1001011011;
    16'b0000000001011000: out_v[329] = 10'b0001001111;
    16'b0001101001010010: out_v[329] = 10'b1011011110;
    16'b0000100000010000: out_v[329] = 10'b1111111000;
    16'b0000001001110000: out_v[329] = 10'b1100010011;
    16'b0001101011010000: out_v[329] = 10'b0110110011;
    16'b0001101001010000: out_v[329] = 10'b1010111001;
    16'b0001100001010000: out_v[329] = 10'b1011000011;
    16'b0000001011010000: out_v[329] = 10'b1110011011;
    16'b0010000000100000: out_v[329] = 10'b0010011010;
    16'b0000101001010000: out_v[329] = 10'b1011101010;
    16'b0000000001100000: out_v[329] = 10'b0110110001;
    16'b0000000000101000: out_v[329] = 10'b1000001100;
    16'b0010000000110000: out_v[329] = 10'b1101011000;
    16'b0000000001101000: out_v[329] = 10'b0100011111;
    16'b0000000000101110: out_v[329] = 10'b0010111000;
    16'b0000000000101010: out_v[329] = 10'b0100100110;
    16'b0000000001001100: out_v[329] = 10'b0000111001;
    16'b0000001000101100: out_v[329] = 10'b0001111101;
    16'b0000000000111010: out_v[329] = 10'b1001111110;
    16'b0000001000111000: out_v[329] = 10'b1001110111;
    16'b0000001000111100: out_v[329] = 10'b0010110110;
    16'b0000000001001000: out_v[329] = 10'b1100101011;
    16'b0000001000101110: out_v[329] = 10'b1100011111;
    16'b0000001000100000: out_v[329] = 10'b0000111101;
    16'b0000001000101000: out_v[329] = 10'b0100110001;
    16'b0000000001101100: out_v[329] = 10'b0110101010;
    16'b0000001000001110: out_v[329] = 10'b0101011001;
    16'b0000001000111110: out_v[329] = 10'b1000111010;
    16'b0000001000001100: out_v[329] = 10'b0101011010;
    16'b0000001000001000: out_v[329] = 10'b0010110001;
    16'b0000001000011100: out_v[329] = 10'b0010110001;
    16'b0000000000111110: out_v[329] = 10'b0010111110;
    16'b0000001000110000: out_v[329] = 10'b0111011011;
    16'b0000000000001110: out_v[329] = 10'b1001110001;
    16'b0000000000010010: out_v[329] = 10'b0110110001;
    16'b0000001001111000: out_v[329] = 10'b1001001010;
    16'b0000000000110010: out_v[329] = 10'b0010110010;
    16'b0000001001100000: out_v[329] = 10'b1110011011;
    16'b0001101001110000: out_v[329] = 10'b0100001000;
    16'b0000101001111000: out_v[329] = 10'b1010111011;
    16'b0001101000110000: out_v[329] = 10'b1011110111;
    16'b0000100000000010: out_v[329] = 10'b0101010010;
    16'b0000100000110010: out_v[329] = 10'b1111010110;
    16'b0000100000010010: out_v[329] = 10'b0011011100;
    16'b0000001001111100: out_v[329] = 10'b0001011110;
    16'b0000000000000010: out_v[329] = 10'b1110101110;
    16'b0000101000110000: out_v[329] = 10'b1101011110;
    16'b0000001001101000: out_v[329] = 10'b1010111111;
    16'b0000000000100010: out_v[329] = 10'b0010100001;
    16'b0001100000000010: out_v[329] = 10'b0010111000;
    16'b0000101000010000: out_v[329] = 10'b1110110111;
    16'b0000000010101000: out_v[329] = 10'b0110100110;
    16'b0010000000001100: out_v[329] = 10'b0011011011;
    16'b0000100010101100: out_v[329] = 10'b0011111000;
    16'b0000000011101100: out_v[329] = 10'b1111111111;
    16'b0001100010101100: out_v[329] = 10'b1010011111;
    16'b0000000010101100: out_v[329] = 10'b1011000000;
    16'b0000000011101000: out_v[329] = 10'b1011001010;
    16'b0000100001101100: out_v[329] = 10'b0100110011;
    16'b0000000010001100: out_v[329] = 10'b0011100110;
    16'b0000000011100000: out_v[329] = 10'b1110111001;
    16'b0000100001001100: out_v[329] = 10'b1001010110;
    16'b0100000000110010: out_v[329] = 10'b0010011110;
    16'b0100000000110000: out_v[329] = 10'b1110111100;
    16'b0000001000110010: out_v[329] = 10'b0110011000;
    16'b0100000000100000: out_v[329] = 10'b1001110011;
    16'b0000010000100000: out_v[329] = 10'b1110001111;
    16'b0100000000100010: out_v[329] = 10'b0101111001;
    16'b0000000000100100: out_v[329] = 10'b1011100000;
    16'b0000010000100010: out_v[329] = 10'b1011010011;
    16'b0000101001110010: out_v[329] = 10'b1011011110;
    16'b0000000001110010: out_v[329] = 10'b0111011010;
    16'b0000101001010010: out_v[329] = 10'b1000011011;
    16'b0000100001110010: out_v[329] = 10'b1111101010;
    16'b0000001001110010: out_v[329] = 10'b0000001001;
    16'b0000001001010010: out_v[329] = 10'b0100001110;
    16'b0000001001100010: out_v[329] = 10'b1111011011;
    16'b0000000001010010: out_v[329] = 10'b1100100110;
    16'b0000001000100010: out_v[329] = 10'b1111000011;
    default: out_v[329] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000100010110001: out_v[330] = 10'b0101000111;
    16'b0001100010110001: out_v[330] = 10'b0110000011;
    16'b1101100011111001: out_v[330] = 10'b1011011110;
    16'b1001100011111000: out_v[330] = 10'b0101101011;
    16'b0000100010110000: out_v[330] = 10'b1101000011;
    16'b0100100011101001: out_v[330] = 10'b1010110101;
    16'b1001100011110001: out_v[330] = 10'b1101011111;
    16'b1001100010110001: out_v[330] = 10'b1010100000;
    16'b1001000011110001: out_v[330] = 10'b0001011011;
    16'b0001100000110001: out_v[330] = 10'b0111110011;
    16'b0000100010011000: out_v[330] = 10'b1101100101;
    16'b0000100011101000: out_v[330] = 10'b1000011101;
    16'b0000100010111000: out_v[330] = 10'b1010101011;
    16'b0001100010110000: out_v[330] = 10'b0110100110;
    16'b1001100010110000: out_v[330] = 10'b0101101010;
    16'b0000100011111000: out_v[330] = 10'b1000111110;
    16'b1101100011101000: out_v[330] = 10'b1111101110;
    16'b1101100011111000: out_v[330] = 10'b1010110010;
    16'b0000100011001000: out_v[330] = 10'b0011000011;
    16'b0100100011111000: out_v[330] = 10'b1110110101;
    16'b1001100011101001: out_v[330] = 10'b0100010111;
    16'b1001100011101000: out_v[330] = 10'b1111010011;
    16'b1001100010010001: out_v[330] = 10'b1101100011;
    16'b0001100010010001: out_v[330] = 10'b1011011110;
    16'b1001100011100000: out_v[330] = 10'b1011001111;
    16'b0100100011101000: out_v[330] = 10'b0101100111;
    16'b1001000010110001: out_v[330] = 10'b1001100010;
    16'b0000100011011000: out_v[330] = 10'b0110111001;
    16'b1101100010110001: out_v[330] = 10'b0000101101;
    16'b0000100010010001: out_v[330] = 10'b1011001010;
    16'b1001000010010001: out_v[330] = 10'b0111010011;
    16'b1001100011110000: out_v[330] = 10'b0011101101;
    16'b0000100000110000: out_v[330] = 10'b1001011100;
    16'b0100100011001000: out_v[330] = 10'b1001011011;
    16'b0000100010111001: out_v[330] = 10'b1101010110;
    16'b1001100011111001: out_v[330] = 10'b0001100110;
    16'b1001100000110001: out_v[330] = 10'b0010110011;
    16'b0001100011111000: out_v[330] = 10'b1110101011;
    16'b0000100011111001: out_v[330] = 10'b0111010011;
    16'b1101100011110001: out_v[330] = 10'b1111011111;
    16'b0100100011111001: out_v[330] = 10'b1011000101;
    16'b0000000010000000: out_v[330] = 10'b0110000110;
    16'b0000000010000001: out_v[330] = 10'b0001001011;
    16'b0000100000000001: out_v[330] = 10'b0010001111;
    16'b0000000000000001: out_v[330] = 10'b0010111010;
    16'b0000100000100001: out_v[330] = 10'b1100001111;
    16'b0000000000100001: out_v[330] = 10'b1001000111;
    16'b0000100010000001: out_v[330] = 10'b0011101000;
    16'b0001000010000000: out_v[330] = 10'b1010010010;
    16'b0001000010000001: out_v[330] = 10'b1100000111;
    16'b0000000000000000: out_v[330] = 10'b0110000111;
    16'b0000100010100001: out_v[330] = 10'b1100010010;
    16'b0000100010000000: out_v[330] = 10'b0000111100;
    16'b1001100010000000: out_v[330] = 10'b0010010100;
    16'b0000000000101001: out_v[330] = 10'b0010101100;
    16'b0000100000000000: out_v[330] = 10'b1000101101;
    16'b1001000010100001: out_v[330] = 10'b1010101110;
    16'b1001000010100000: out_v[330] = 10'b0010011111;
    16'b0000100010001000: out_v[330] = 10'b0100001101;
    16'b1001000000010000: out_v[330] = 10'b1011101101;
    16'b1001000010010000: out_v[330] = 10'b0100000110;
    16'b1001000000000000: out_v[330] = 10'b1011110110;
    16'b0000000010100000: out_v[330] = 10'b0110110101;
    16'b1001000010000000: out_v[330] = 10'b1111001010;
    16'b1001100010010000: out_v[330] = 10'b0001011100;
    16'b0000000000010000: out_v[330] = 10'b0110101101;
    16'b0001000010010000: out_v[330] = 10'b0010100110;
    16'b0000100010010000: out_v[330] = 10'b0110000100;
    16'b0000000010010000: out_v[330] = 10'b1010000100;
    16'b0001000010100000: out_v[330] = 10'b1111010101;
    16'b0000100010101000: out_v[330] = 10'b1010001110;
    16'b1001000010001000: out_v[330] = 10'b1010100111;
    16'b1001000010110000: out_v[330] = 10'b0111000110;
    16'b0001100010000000: out_v[330] = 10'b0010011011;
    16'b0001000010001000: out_v[330] = 10'b1101111100;
    16'b1001000010101000: out_v[330] = 10'b1010010110;
    16'b0001100010101000: out_v[330] = 10'b1010011101;
    16'b1001000000100000: out_v[330] = 10'b0111110001;
    16'b0000000010101000: out_v[330] = 10'b0110010011;
    16'b0001000010101000: out_v[330] = 10'b1011010111;
    16'b0001100010100000: out_v[330] = 10'b1011011111;
    16'b0000100010101001: out_v[330] = 10'b0011110000;
    16'b0000100010100000: out_v[330] = 10'b1100100010;
    16'b0000100010001001: out_v[330] = 10'b1011010011;
    16'b0000000010100001: out_v[330] = 10'b0110101000;
    16'b0000000010010001: out_v[330] = 10'b0011011000;
    16'b0000000010001000: out_v[330] = 10'b1110100001;
    16'b0001100010001000: out_v[330] = 10'b1100001011;
    16'b0000000000010001: out_v[330] = 10'b0100111001;
    16'b1000000000010000: out_v[330] = 10'b1011100110;
    16'b1001100010100000: out_v[330] = 10'b0010111011;
    16'b1001100010100001: out_v[330] = 10'b1011011110;
    16'b0000100000001000: out_v[330] = 10'b0100110110;
    16'b0000100000010001: out_v[330] = 10'b0100001011;
    16'b0000100000010000: out_v[330] = 10'b0010111101;
    16'b1001100010000001: out_v[330] = 10'b0011111001;
    16'b0000100010011001: out_v[330] = 10'b0110010111;
    16'b0000100000111001: out_v[330] = 10'b0010101111;
    16'b0001100010010000: out_v[330] = 10'b0111111010;
    16'b0000100000100000: out_v[330] = 10'b0111110001;
    16'b0001100010000001: out_v[330] = 10'b1100010000;
    16'b0000100000001001: out_v[330] = 10'b1101000001;
    16'b1001000010000001: out_v[330] = 10'b0110111000;
    16'b0001100000000001: out_v[330] = 10'b0011110011;
    16'b0001100000010001: out_v[330] = 10'b1101001101;
    16'b0000100000101000: out_v[330] = 10'b0011101011;
    16'b0000100000101001: out_v[330] = 10'b0111111100;
    16'b0000100000011001: out_v[330] = 10'b0001010010;
    16'b0001100010100001: out_v[330] = 10'b1101011100;
    16'b1001100010101000: out_v[330] = 10'b1000011110;
    16'b0000100000110001: out_v[330] = 10'b0111011000;
    16'b0000000000111000: out_v[330] = 10'b0011110110;
    16'b0000100001110000: out_v[330] = 10'b1000011101;
    16'b0000000000011000: out_v[330] = 10'b0101110101;
    16'b0000000000110000: out_v[330] = 10'b0101011011;
    16'b0000000001001000: out_v[330] = 10'b1001011000;
    16'b0000000010110000: out_v[330] = 10'b1001001011;
    16'b0000100001111000: out_v[330] = 10'b1000101110;
    16'b0000100000011000: out_v[330] = 10'b1011000011;
    16'b0000100001011000: out_v[330] = 10'b0010110001;
    16'b0000000001111000: out_v[330] = 10'b0110111100;
    16'b0000000001011000: out_v[330] = 10'b1101000111;
    16'b0000000010110001: out_v[330] = 10'b1111101110;
    16'b0000100000111000: out_v[330] = 10'b1011000000;
    16'b0000100001001000: out_v[330] = 10'b0011110100;
    16'b0000000001010100: out_v[330] = 10'b0100110010;
    16'b0000000001110000: out_v[330] = 10'b0101010111;
    16'b0000100001110001: out_v[330] = 10'b0100011000;
    16'b0000000000100000: out_v[330] = 10'b0001111011;
    16'b0000000000011001: out_v[330] = 10'b1001011101;
    16'b0000000001010000: out_v[330] = 10'b0001101111;
    16'b0000000000110001: out_v[330] = 10'b1010101010;
    16'b0000000011110000: out_v[330] = 10'b1011000110;
    16'b0001000010010001: out_v[330] = 10'b1101000011;
    16'b0001000010110001: out_v[330] = 10'b0011101110;
    16'b0001100000110000: out_v[330] = 10'b0101110110;
    16'b0010100000110001: out_v[330] = 10'b0010110111;
    16'b0010100010110001: out_v[330] = 10'b1000111111;
    16'b0100000001011000: out_v[330] = 10'b1110111001;
    16'b0000000010111000: out_v[330] = 10'b1101100011;
    16'b0100000001001000: out_v[330] = 10'b0101101010;
    16'b0100000010110000: out_v[330] = 10'b1010111100;
    16'b0000000000101101: out_v[330] = 10'b1101110110;
    16'b0000000000101000: out_v[330] = 10'b0111011010;
    16'b0000100001100001: out_v[330] = 10'b1011100110;
    16'b0000100001101001: out_v[330] = 10'b0011101111;
    16'b0000000010101001: out_v[330] = 10'b1010100010;
    16'b0000000001101001: out_v[330] = 10'b1111000110;
    16'b0000100000101100: out_v[330] = 10'b0111101011;
    16'b0000100000101101: out_v[330] = 10'b1100101011;
    16'b0000000000111001: out_v[330] = 10'b1111011100;
    16'b0000100000101111: out_v[330] = 10'b0011010011;
    16'b0000100001111001: out_v[330] = 10'b0110000000;
    16'b0000100001101101: out_v[330] = 10'b0011101010;
    16'b0000000000101111: out_v[330] = 10'b0110010110;
    16'b0000100001101000: out_v[330] = 10'b0110100010;
    16'b0000000001101101: out_v[330] = 10'b0011000101;
    16'b0001100000100000: out_v[330] = 10'b1100100111;
    16'b0001100000100001: out_v[330] = 10'b1101100010;
    16'b0000000001101000: out_v[330] = 10'b1000101000;
    16'b0000000001100000: out_v[330] = 10'b1001110011;
    16'b0000000001111001: out_v[330] = 10'b1001100010;
    16'b0000100001100000: out_v[330] = 10'b1000011101;
    default: out_v[330] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001100001001000: out_v[331] = 10'b1011011010;
    16'b0101100000011100: out_v[331] = 10'b1111011111;
    16'b0000100001000100: out_v[331] = 10'b0000110101;
    16'b0000000001000000: out_v[331] = 10'b1000111100;
    16'b0000100001001000: out_v[331] = 10'b1011110000;
    16'b0000100000011100: out_v[331] = 10'b0101010001;
    16'b0000100000001100: out_v[331] = 10'b1100000010;
    16'b0000100001010100: out_v[331] = 10'b0100000001;
    16'b0000100001010000: out_v[331] = 10'b0110110110;
    16'b0000000000000000: out_v[331] = 10'b0101101101;
    16'b0000100001001100: out_v[331] = 10'b0110111101;
    16'b0101100001000000: out_v[331] = 10'b0011011101;
    16'b0101000001000000: out_v[331] = 10'b1100110101;
    16'b0101000001001000: out_v[331] = 10'b1001001010;
    16'b0101000000000000: out_v[331] = 10'b0100111100;
    16'b0000100000000100: out_v[331] = 10'b1101010110;
    16'b0000100000000000: out_v[331] = 10'b0111001110;
    16'b0000100000001000: out_v[331] = 10'b1100111001;
    16'b0000000001001000: out_v[331] = 10'b1001011110;
    16'b0000100001000000: out_v[331] = 10'b1001100111;
    16'b0000100000010100: out_v[331] = 10'b0001010011;
    16'b0101100001011100: out_v[331] = 10'b0000010001;
    16'b0001000001001000: out_v[331] = 10'b1111001001;
    16'b0000100001011100: out_v[331] = 10'b0000011011;
    16'b0101100001010100: out_v[331] = 10'b0000111001;
    16'b0101100001001000: out_v[331] = 10'b1110001010;
    16'b0101100001001100: out_v[331] = 10'b1101101110;
    16'b0101100001000100: out_v[331] = 10'b0101011001;
    16'b0001000001000000: out_v[331] = 10'b1101101001;
    16'b0000100001011000: out_v[331] = 10'b0011101011;
    16'b0000100000011000: out_v[331] = 10'b1000000101;
    16'b0000100001001001: out_v[331] = 10'b1011001011;
    16'b0000000000001000: out_v[331] = 10'b0110011110;
    16'b0100000000001000: out_v[331] = 10'b0000110011;
    16'b0100000000000000: out_v[331] = 10'b0110110011;
    16'b0001000000001000: out_v[331] = 10'b0010100010;
    16'b0101000000001000: out_v[331] = 10'b1010001110;
    16'b0100000001001000: out_v[331] = 10'b1110000110;
    16'b0000000000000001: out_v[331] = 10'b1111011010;
    16'b0000000001000010: out_v[331] = 10'b0101110110;
    16'b0000000000001010: out_v[331] = 10'b0001100110;
    16'b0000000000100000: out_v[331] = 10'b1110010100;
    16'b0000000001010000: out_v[331] = 10'b1010100111;
    16'b0000000000000010: out_v[331] = 10'b1010000101;
    16'b0000000000010000: out_v[331] = 10'b0110100100;
    16'b0000000000011000: out_v[331] = 10'b1100001110;
    16'b0000000000110000: out_v[331] = 10'b1100010101;
    16'b0000000100000000: out_v[331] = 10'b1001000000;
    16'b0000000000101000: out_v[331] = 10'b0110110110;
    16'b0000000000111000: out_v[331] = 10'b0100101111;
    16'b0000000101000000: out_v[331] = 10'b1010010100;
    16'b0001000000000000: out_v[331] = 10'b0110010001;
    16'b0101100000000100: out_v[331] = 10'b0001110001;
    16'b0001100000000000: out_v[331] = 10'b0010110101;
    16'b0001100000000100: out_v[331] = 10'b1101010011;
    16'b0000110000000100: out_v[331] = 10'b1000010110;
    16'b0000100000000101: out_v[331] = 10'b0010110011;
    16'b0100100000000100: out_v[331] = 10'b1100110111;
    16'b0001100001000000: out_v[331] = 10'b1100101010;
    16'b0100100000000000: out_v[331] = 10'b0110110111;
    16'b0100000001000000: out_v[331] = 10'b0111010001;
    16'b0100100001000100: out_v[331] = 10'b1111100010;
    16'b0000110000000000: out_v[331] = 10'b0111110110;
    16'b0100100001000000: out_v[331] = 10'b1000100000;
    16'b0100110000000100: out_v[331] = 10'b0100111001;
    16'b0000100000010000: out_v[331] = 10'b1001001000;
    16'b0000100000000001: out_v[331] = 10'b1010111010;
    16'b0101100000000000: out_v[331] = 10'b0001011110;
    16'b0100100000001000: out_v[331] = 10'b0111100110;
    16'b0101100000001000: out_v[331] = 10'b0110101111;
    16'b0000000001000001: out_v[331] = 10'b1000100000;
    16'b0101100000001100: out_v[331] = 10'b0011100111;
    16'b0000000001001001: out_v[331] = 10'b1001100011;
    16'b0000100000110100: out_v[331] = 10'b0111110011;
    16'b0000100100010100: out_v[331] = 10'b1001011000;
    16'b0000100100010000: out_v[331] = 10'b1100101011;
    16'b0000100100000000: out_v[331] = 10'b0111001010;
    16'b0000000100010000: out_v[331] = 10'b1111100000;
    16'b0100100000001100: out_v[331] = 10'b1111100001;
    16'b0000010000001000: out_v[331] = 10'b1001101001;
    16'b0100010000001000: out_v[331] = 10'b0110110101;
    16'b0100010000000000: out_v[331] = 10'b1100001101;
    16'b0001100000001000: out_v[331] = 10'b0011101011;
    16'b0001100000001100: out_v[331] = 10'b1101101110;
    16'b0000010000000000: out_v[331] = 10'b1111001001;
    16'b0101000000001100: out_v[331] = 10'b0011011101;
    16'b0100000010001000: out_v[331] = 10'b1101100101;
    16'b0000110000001100: out_v[331] = 10'b1101001001;
    16'b0100010010001000: out_v[331] = 10'b1001110111;
    16'b0100110010001100: out_v[331] = 10'b1101000111;
    16'b0100000010000000: out_v[331] = 10'b1101001110;
    16'b0101000010001000: out_v[331] = 10'b0001111111;
    16'b0001000000001100: out_v[331] = 10'b1100111111;
    16'b0100100010001100: out_v[331] = 10'b1111011010;
    16'b0001100001000100: out_v[331] = 10'b1111000110;
    16'b0000110000001000: out_v[331] = 10'b1001100111;
    16'b0100110000000000: out_v[331] = 10'b1110101010;
    16'b0100100010000000: out_v[331] = 10'b1010001111;
    16'b0100100010001000: out_v[331] = 10'b1111100111;
    16'b0100110000001100: out_v[331] = 10'b0000111110;
    16'b0100110000001000: out_v[331] = 10'b1011101110;
    default: out_v[331] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001000011100010: out_v[332] = 10'b1001000101;
    16'b0001000111100000: out_v[332] = 10'b0011101110;
    16'b0001000001100010: out_v[332] = 10'b0100010001;
    16'b0000000011100010: out_v[332] = 10'b1101010011;
    16'b0000000011100000: out_v[332] = 10'b0101010011;
    16'b0001000010001000: out_v[332] = 10'b1000011111;
    16'b0000000010001000: out_v[332] = 10'b1001010011;
    16'b0000000011101000: out_v[332] = 10'b0000011101;
    16'b0000000011101010: out_v[332] = 10'b0101001111;
    16'b0001000011100000: out_v[332] = 10'b0101010101;
    16'b1001000001100010: out_v[332] = 10'b0110110111;
    16'b0001000001100000: out_v[332] = 10'b1000101011;
    16'b0001000011101010: out_v[332] = 10'b1110000110;
    16'b0001000010100010: out_v[332] = 10'b1100100110;
    16'b0000000000001000: out_v[332] = 10'b1011000011;
    16'b0001000010100000: out_v[332] = 10'b0101101010;
    16'b0000000111100000: out_v[332] = 10'b0011100001;
    16'b0001000011101000: out_v[332] = 10'b1110001101;
    16'b0000000111100010: out_v[332] = 10'b0000001111;
    16'b0000000111101000: out_v[332] = 10'b0011001010;
    16'b0001000010000010: out_v[332] = 10'b0110110000;
    16'b0000000001100010: out_v[332] = 10'b0010110110;
    16'b0000000010101000: out_v[332] = 10'b1100111000;
    16'b1001000011100010: out_v[332] = 10'b0110010011;
    16'b0001000000100010: out_v[332] = 10'b0101001100;
    16'b0001000000100000: out_v[332] = 10'b0011001011;
    16'b1001010000101100: out_v[332] = 10'b1100110010;
    16'b0001000000000010: out_v[332] = 10'b1011101000;
    16'b0001000010101000: out_v[332] = 10'b0111110110;
    16'b1001000000101000: out_v[332] = 10'b0011100110;
    16'b0001000000001000: out_v[332] = 10'b1001011110;
    16'b1001010000001100: out_v[332] = 10'b1101010011;
    16'b1001000000001000: out_v[332] = 10'b1111000011;
    16'b0001000111100010: out_v[332] = 10'b1111011010;
    16'b0000000000000000: out_v[332] = 10'b1011011001;
    16'b0001000000000000: out_v[332] = 10'b0010000111;
    16'b0000000010000000: out_v[332] = 10'b1101100010;
    16'b0001000010000000: out_v[332] = 10'b1110100111;
    16'b0010000010000000: out_v[332] = 10'b1011011011;
    16'b0000000000000010: out_v[332] = 10'b1111101010;
    16'b0000000100000010: out_v[332] = 10'b0111000111;
    16'b0000000100000000: out_v[332] = 10'b0110100010;
    16'b0110000000000000: out_v[332] = 10'b1100100100;
    16'b0110000010000000: out_v[332] = 10'b1010001111;
    16'b0110000001100010: out_v[332] = 10'b0111010110;
    16'b0111000000000000: out_v[332] = 10'b0100110011;
    16'b1000000000000000: out_v[332] = 10'b0111110001;
    16'b0000000000100000: out_v[332] = 10'b1011101111;
    16'b0000000000100010: out_v[332] = 10'b1100100110;
    16'b1001010000000100: out_v[332] = 10'b1101110110;
    16'b0110000000100010: out_v[332] = 10'b1001100101;
    16'b1000010000000100: out_v[332] = 10'b0101110101;
    16'b0010000000100010: out_v[332] = 10'b0011001001;
    16'b0110000000000010: out_v[332] = 10'b1001100111;
    16'b0000000001100000: out_v[332] = 10'b0111011000;
    16'b1001010000000000: out_v[332] = 10'b1101010100;
    16'b0000000010100010: out_v[332] = 10'b1110000111;
    16'b1000010000000110: out_v[332] = 10'b0010111000;
    16'b0000000000101010: out_v[332] = 10'b1101111110;
    16'b0000000001101010: out_v[332] = 10'b0011100111;
    16'b1000010000100110: out_v[332] = 10'b1000101111;
    16'b0000000010100000: out_v[332] = 10'b1110110100;
    16'b0010000000000010: out_v[332] = 10'b1111111111;
    16'b1000000000000010: out_v[332] = 10'b0010111100;
    16'b1001010000000010: out_v[332] = 10'b0001110010;
    16'b1000000000100010: out_v[332] = 10'b1010110010;
    16'b0111000000000010: out_v[332] = 10'b1000001110;
    16'b1001010000000110: out_v[332] = 10'b0001001100;
    16'b0010000000100000: out_v[332] = 10'b1100101011;
    16'b1000010000100010: out_v[332] = 10'b1001110111;
    16'b0010000000000000: out_v[332] = 10'b1001110101;
    16'b1000010010000100: out_v[332] = 10'b0010011110;
    16'b0110000000100000: out_v[332] = 10'b0111000110;
    16'b0110000010100000: out_v[332] = 10'b0100011111;
    16'b1000010000000010: out_v[332] = 10'b0111011011;
    16'b0000000010000010: out_v[332] = 10'b0011011100;
    16'b1000010000000000: out_v[332] = 10'b0011010011;
    16'b0000000100100010: out_v[332] = 10'b0010011110;
    16'b1110010000100010: out_v[332] = 10'b0010011000;
    16'b1001010010000100: out_v[332] = 10'b1011001010;
    16'b0001000001000010: out_v[332] = 10'b1100010001;
    16'b1001010010000000: out_v[332] = 10'b1111011111;
    16'b0111000001000000: out_v[332] = 10'b1110101010;
    16'b1001000000000000: out_v[332] = 10'b0000111101;
    16'b0001000001000000: out_v[332] = 10'b0110110101;
    16'b0011000010000010: out_v[332] = 10'b0110011001;
    16'b1001010010000110: out_v[332] = 10'b1110001110;
    16'b1001000010000000: out_v[332] = 10'b0001001100;
    16'b0011000010000000: out_v[332] = 10'b0111001010;
    16'b0001000011000010: out_v[332] = 10'b1100101000;
    16'b0110000010000010: out_v[332] = 10'b1011011010;
    16'b0111000010000000: out_v[332] = 10'b1111011011;
    16'b1001010010000010: out_v[332] = 10'b1111110110;
    16'b0011000000000000: out_v[332] = 10'b0011111100;
    16'b0111000011000000: out_v[332] = 10'b0001001111;
    16'b1001010011000100: out_v[332] = 10'b1011111110;
    16'b1001000000000010: out_v[332] = 10'b1001010010;
    16'b0111000010000010: out_v[332] = 10'b1101011111;
    16'b1001010001000000: out_v[332] = 10'b0011111100;
    16'b0001000011000000: out_v[332] = 10'b1001110011;
    16'b1000000001100010: out_v[332] = 10'b0010111101;
    16'b1000000001100000: out_v[332] = 10'b0011110111;
    16'b0000000001000000: out_v[332] = 10'b1100111000;
    16'b1000010001100010: out_v[332] = 10'b0110110010;
    16'b0000000101100010: out_v[332] = 10'b1100111011;
    16'b1000010001000110: out_v[332] = 10'b1101001000;
    16'b0001000101101010: out_v[332] = 10'b1011100111;
    16'b1000010001101110: out_v[332] = 10'b1100011111;
    16'b1000010001100110: out_v[332] = 10'b1111001110;
    16'b1000010001000000: out_v[332] = 10'b1000100010;
    16'b1000010001000010: out_v[332] = 10'b0011010000;
    16'b0000000001000010: out_v[332] = 10'b1001111011;
    16'b1000010001100000: out_v[332] = 10'b0000111111;
    16'b0000000111101010: out_v[332] = 10'b0010111111;
    16'b1000010000101110: out_v[332] = 10'b1101110000;
    16'b1000000001101010: out_v[332] = 10'b1011011111;
    16'b1000000001000000: out_v[332] = 10'b0110010001;
    16'b0000000011000010: out_v[332] = 10'b0101110100;
    16'b0000000101101010: out_v[332] = 10'b0011101110;
    16'b0001000101100010: out_v[332] = 10'b0110111110;
    16'b1000000001000010: out_v[332] = 10'b1100000111;
    16'b0001000111101010: out_v[332] = 10'b1010000110;
    16'b0000000011000000: out_v[332] = 10'b1101010110;
    16'b0001000110000000: out_v[332] = 10'b1010110110;
    16'b0001000111000000: out_v[332] = 10'b1000011111;
    16'b0000000111000000: out_v[332] = 10'b1110100100;
    16'b0001000101000000: out_v[332] = 10'b1101011010;
    16'b0000000110000000: out_v[332] = 10'b0110100101;
    16'b0001000100000000: out_v[332] = 10'b0101001100;
    16'b0001000101100000: out_v[332] = 10'b0001111111;
    16'b1001000001000000: out_v[332] = 10'b0011110010;
    16'b0000000110100000: out_v[332] = 10'b0010111010;
    16'b1110010001100110: out_v[332] = 10'b1101001011;
    16'b1110010001100010: out_v[332] = 10'b1010001001;
    16'b1010000001100010: out_v[332] = 10'b1111000110;
    16'b0010000001100010: out_v[332] = 10'b1010111001;
    16'b1110000001100010: out_v[332] = 10'b1111101011;
    16'b1110010000100110: out_v[332] = 10'b1101001001;
    16'b0000000010000110: out_v[332] = 10'b0000011101;
    16'b1000010010000110: out_v[332] = 10'b1011011000;
    16'b1000010010000010: out_v[332] = 10'b0110101110;
    16'b1001000010000010: out_v[332] = 10'b0111001010;
    16'b1000010010000000: out_v[332] = 10'b1100011100;
    16'b1000000010000010: out_v[332] = 10'b1000101111;
    16'b0001000010000110: out_v[332] = 10'b0011111000;
    16'b0001000110100010: out_v[332] = 10'b1101001111;
    16'b0001000110000010: out_v[332] = 10'b0010110110;
    16'b1001010001000110: out_v[332] = 10'b1101000010;
    16'b0001000100000010: out_v[332] = 10'b1001001111;
    16'b1001010001100110: out_v[332] = 10'b1110001110;
    16'b0000000110100010: out_v[332] = 10'b1110100101;
    16'b0000000110000010: out_v[332] = 10'b1101100110;
    16'b0000000010101010: out_v[332] = 10'b1100101010;
    16'b1001000001000010: out_v[332] = 10'b1000100111;
    default: out_v[332] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010101000000011: out_v[333] = 10'b0010001011;
    16'b0010101000001011: out_v[333] = 10'b0001110001;
    16'b0000101000000001: out_v[333] = 10'b0000100101;
    16'b0000100000000011: out_v[333] = 10'b1011110100;
    16'b0000100000000010: out_v[333] = 10'b1011100101;
    16'b0000101000000011: out_v[333] = 10'b1000101011;
    16'b0000101000000010: out_v[333] = 10'b1101110110;
    16'b0000101000001011: out_v[333] = 10'b1000010111;
    16'b0010100000000010: out_v[333] = 10'b0101111111;
    16'b0100100000000001: out_v[333] = 10'b0100111011;
    16'b0010100000000011: out_v[333] = 10'b1110110110;
    16'b0000100000000001: out_v[333] = 10'b0101000101;
    16'b0110101000000011: out_v[333] = 10'b0000011000;
    16'b0100101000000011: out_v[333] = 10'b1010100010;
    16'b0000101000001001: out_v[333] = 10'b1011110001;
    16'b0100100000000011: out_v[333] = 10'b1110101001;
    16'b0000001000000010: out_v[333] = 10'b0101000010;
    16'b0000000000000010: out_v[333] = 10'b0111110101;
    16'b0000100000000000: out_v[333] = 10'b1010001101;
    16'b0100101000000001: out_v[333] = 10'b0010011010;
    16'b0010101000000010: out_v[333] = 10'b0101011000;
    16'b0100001000000001: out_v[333] = 10'b0100011011;
    16'b0010000000000010: out_v[333] = 10'b0110010100;
    16'b0000001000001010: out_v[333] = 10'b0110100001;
    16'b0010100000000001: out_v[333] = 10'b0011110000;
    16'b0100000000000001: out_v[333] = 10'b1100110011;
    16'b0000101000001010: out_v[333] = 10'b0111001111;
    16'b0000100000001011: out_v[333] = 10'b0010101111;
    16'b0010101000000001: out_v[333] = 10'b0111100111;
    16'b0000000000000000: out_v[333] = 10'b1100010000;
    16'b0010000000000000: out_v[333] = 10'b1000011000;
    16'b0000001000000000: out_v[333] = 10'b1001001101;
    16'b0100000000000010: out_v[333] = 10'b1010011110;
    16'b0100000000000100: out_v[333] = 10'b1001100101;
    16'b0100010000000000: out_v[333] = 10'b1100100100;
    16'b0100000000000000: out_v[333] = 10'b1001110110;
    16'b0000101000000000: out_v[333] = 10'b0110001010;
    16'b0000111000000000: out_v[333] = 10'b1010001001;
    16'b0000010000000000: out_v[333] = 10'b1101100110;
    16'b0100100000000100: out_v[333] = 10'b1011000010;
    16'b0100010000000100: out_v[333] = 10'b1111100101;
    16'b0100101000000100: out_v[333] = 10'b1111100101;
    16'b0100101000000000: out_v[333] = 10'b1111000101;
    16'b0100001000000000: out_v[333] = 10'b0101110011;
    16'b0000000000000001: out_v[333] = 10'b1111010011;
    16'b0000111000000001: out_v[333] = 10'b0110110111;
    16'b0000110000000000: out_v[333] = 10'b1101010111;
    16'b0001101000000000: out_v[333] = 10'b0110010111;
    16'b0101001000000000: out_v[333] = 10'b0101010110;
    16'b0100001000000100: out_v[333] = 10'b1011000111;
    16'b0000110000000001: out_v[333] = 10'b1011100101;
    16'b0001001000000000: out_v[333] = 10'b1011000111;
    16'b0100100000000000: out_v[333] = 10'b0101010000;
    16'b0000001000000001: out_v[333] = 10'b1000100111;
    16'b0000000000000011: out_v[333] = 10'b0010111101;
    16'b0001101000000001: out_v[333] = 10'b1010111101;
    16'b0100001000000010: out_v[333] = 10'b0011110110;
    16'b0010100000000000: out_v[333] = 10'b0110110011;
    16'b0110100000000000: out_v[333] = 10'b0011011111;
    16'b0010101000000000: out_v[333] = 10'b1011001110;
    16'b0100100000000101: out_v[333] = 10'b0111111001;
    16'b0110101000000001: out_v[333] = 10'b0111011111;
    16'b0100100000000111: out_v[333] = 10'b1111001100;
    16'b0110100000000001: out_v[333] = 10'b1011110011;
    16'b0110100000000011: out_v[333] = 10'b1000010110;
    16'b0100100000000010: out_v[333] = 10'b0101001001;
    16'b0110100000000101: out_v[333] = 10'b1001100101;
    16'b0000110000000011: out_v[333] = 10'b1110011000;
    16'b0000111000000011: out_v[333] = 10'b1000001011;
    16'b0010001000000000: out_v[333] = 10'b0110001001;
    16'b0100100000000110: out_v[333] = 10'b0111011001;
    16'b0000100000000101: out_v[333] = 10'b1000011011;
    16'b0000000000001010: out_v[333] = 10'b1110101110;
    16'b0010001000000010: out_v[333] = 10'b1111110010;
    16'b0000001000010010: out_v[333] = 10'b1110001000;
    16'b0110100000000010: out_v[333] = 10'b1000011010;
    16'b0000000000010010: out_v[333] = 10'b0010111101;
    16'b0100000000000101: out_v[333] = 10'b0110001010;
    16'b0010000000010010: out_v[333] = 10'b1100000011;
    16'b0001100000000010: out_v[333] = 10'b1101000111;
    16'b0001100000000011: out_v[333] = 10'b1001000010;
    16'b0001000000000010: out_v[333] = 10'b0110101000;
    16'b0001000000000000: out_v[333] = 10'b1011100011;
    16'b0001101000000011: out_v[333] = 10'b1011011010;
    16'b0000100000001001: out_v[333] = 10'b0011001111;
    16'b0000110000100001: out_v[333] = 10'b1001001010;
    16'b0001100000000000: out_v[333] = 10'b1001001011;
    16'b0001101000000010: out_v[333] = 10'b0011011011;
    16'b0010000100000010: out_v[333] = 10'b0110101001;
    16'b0000000100000010: out_v[333] = 10'b1111001101;
    16'b0010000100000000: out_v[333] = 10'b1001111111;
    16'b0010001000001010: out_v[333] = 10'b0100110000;
    16'b0010000000001010: out_v[333] = 10'b1001100110;
    default: out_v[333] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1000001000000000: out_v[334] = 10'b0010101011;
    16'b1000001000001000: out_v[334] = 10'b1110000001;
    16'b1000001000001010: out_v[334] = 10'b0010010011;
    16'b0000001000011010: out_v[334] = 10'b0111000111;
    16'b0000000000000010: out_v[334] = 10'b1000110000;
    16'b1000001000011000: out_v[334] = 10'b1101000111;
    16'b0000000000000000: out_v[334] = 10'b0001011000;
    16'b0000000000001010: out_v[334] = 10'b0111010100;
    16'b0000001000000010: out_v[334] = 10'b0110010010;
    16'b0000001000000000: out_v[334] = 10'b1100111100;
    16'b0000001000001010: out_v[334] = 10'b0101001010;
    16'b0000000000001000: out_v[334] = 10'b0101100001;
    16'b0000001000001000: out_v[334] = 10'b0111111101;
    16'b1000000000000000: out_v[334] = 10'b0100010010;
    16'b1000000000001010: out_v[334] = 10'b0110011011;
    16'b1000011000001010: out_v[334] = 10'b1100000111;
    16'b0000011000000010: out_v[334] = 10'b1000001100;
    16'b1000000000001000: out_v[334] = 10'b0011110001;
    16'b1000001001001000: out_v[334] = 10'b0011010101;
    16'b0000010000001010: out_v[334] = 10'b0100010111;
    16'b1000001001011000: out_v[334] = 10'b1000111011;
    16'b0000001000011000: out_v[334] = 10'b0110100011;
    16'b0010011000001010: out_v[334] = 10'b1111111011;
    16'b1000001000000010: out_v[334] = 10'b0010101011;
    16'b0000011000001010: out_v[334] = 10'b1100011110;
    16'b1000001000011010: out_v[334] = 10'b1100110101;
    16'b1010011000001010: out_v[334] = 10'b0010010101;
    16'b1000000000000010: out_v[334] = 10'b1000100110;
    16'b1000010000000000: out_v[334] = 10'b1011011100;
    16'b0000011000000000: out_v[334] = 10'b0100111100;
    16'b1010001000000000: out_v[334] = 10'b0011101110;
    16'b0010000000000000: out_v[334] = 10'b0001110100;
    16'b0000010000000010: out_v[334] = 10'b0001110110;
    16'b0010001000000000: out_v[334] = 10'b1001010010;
    16'b1010001000000010: out_v[334] = 10'b0011110100;
    16'b0000000000011000: out_v[334] = 10'b0010000101;
    16'b0000010000000000: out_v[334] = 10'b0101010111;
    16'b0010001000000010: out_v[334] = 10'b0100100100;
    16'b0000001001000000: out_v[334] = 10'b1100000010;
    16'b0011001000000010: out_v[334] = 10'b1001110100;
    16'b0000000001000010: out_v[334] = 10'b1001111011;
    16'b0010000000000010: out_v[334] = 10'b1111011000;
    16'b0000000001000000: out_v[334] = 10'b0011001111;
    16'b0011001000000000: out_v[334] = 10'b1000100011;
    16'b1000001001000000: out_v[334] = 10'b1010101100;
    16'b0000000000010000: out_v[334] = 10'b1110001111;
    16'b0010011000000010: out_v[334] = 10'b1111001011;
    16'b1000011000000000: out_v[334] = 10'b1011100111;
    16'b0000001000010000: out_v[334] = 10'b0010001100;
    16'b1000011000000010: out_v[334] = 10'b1100101100;
    16'b0000001001000010: out_v[334] = 10'b0011001011;
    16'b1000010000000010: out_v[334] = 10'b1000101010;
    16'b0000011000100000: out_v[334] = 10'b0111110011;
    16'b0000000000001110: out_v[334] = 10'b0111110011;
    16'b0000000000001100: out_v[334] = 10'b0101010011;
    16'b0000000000000110: out_v[334] = 10'b0111001011;
    16'b1000001000101000: out_v[334] = 10'b1000011011;
    16'b1000101000000000: out_v[334] = 10'b1010001110;
    16'b0000000000101000: out_v[334] = 10'b0111001110;
    16'b1000001000100000: out_v[334] = 10'b1001011111;
    16'b0000011000100010: out_v[334] = 10'b1001100110;
    default: out_v[334] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001100010101100: out_v[335] = 10'b0001011000;
    16'b0111000111111101: out_v[335] = 10'b0111001110;
    16'b0000100010101100: out_v[335] = 10'b0110101001;
    16'b0001100010101000: out_v[335] = 10'b0110011011;
    16'b0001100010100100: out_v[335] = 10'b0000101001;
    16'b0011100010101100: out_v[335] = 10'b0111101110;
    16'b0011100110111000: out_v[335] = 10'b1110101011;
    16'b0001100011101100: out_v[335] = 10'b1100010111;
    16'b0000100010101000: out_v[335] = 10'b0010100011;
    16'b0111000101111001: out_v[335] = 10'b1100110010;
    16'b0111000111101101: out_v[335] = 10'b0111010011;
    16'b0011000111111101: out_v[335] = 10'b0110110111;
    16'b0011000110101100: out_v[335] = 10'b1011110011;
    16'b0111001111011101: out_v[335] = 10'b0101111110;
    16'b0111000111011101: out_v[335] = 10'b0011010101;
    16'b0011100110111100: out_v[335] = 10'b0100100110;
    16'b0011000111111100: out_v[335] = 10'b0111111110;
    16'b0011100111101100: out_v[335] = 10'b0010111011;
    16'b0011100110001000: out_v[335] = 10'b1110111111;
    16'b0110000111111101: out_v[335] = 10'b1101011111;
    16'b0011100110101000: out_v[335] = 10'b1100010110;
    16'b0011100110101100: out_v[335] = 10'b0100001001;
    16'b0111000111111001: out_v[335] = 10'b0010101101;
    16'b0111100111111101: out_v[335] = 10'b1000011011;
    16'b0011100111111100: out_v[335] = 10'b1111001110;
    16'b0001100010001000: out_v[335] = 10'b1000101111;
    16'b0000100010001100: out_v[335] = 10'b0111111001;
    16'b0011000110111100: out_v[335] = 10'b0011101110;
    16'b0011100111111101: out_v[335] = 10'b1011111111;
    16'b0001100010000100: out_v[335] = 10'b1110100111;
    16'b0000100010100100: out_v[335] = 10'b0001100110;
    16'b0011000111101100: out_v[335] = 10'b1101111010;
    16'b0011000111101101: out_v[335] = 10'b1101111101;
    16'b0001000011101100: out_v[335] = 10'b0101001001;
    16'b0111001111111101: out_v[335] = 10'b0101010111;
    16'b0011100110110100: out_v[335] = 10'b1000110001;
    16'b0001100010001100: out_v[335] = 10'b1110001010;
    16'b0001000010000000: out_v[335] = 10'b0110101011;
    16'b0000000000000100: out_v[335] = 10'b1001011111;
    16'b0000000000000000: out_v[335] = 10'b1000000111;
    16'b0000000010000100: out_v[335] = 10'b0100100001;
    16'b0001000000000000: out_v[335] = 10'b0110000011;
    16'b0000000010000000: out_v[335] = 10'b1000111011;
    16'b0000000010001000: out_v[335] = 10'b0110001000;
    16'b0001000010000100: out_v[335] = 10'b0001111111;
    16'b0001000000000100: out_v[335] = 10'b0111110000;
    16'b0001000010001000: out_v[335] = 10'b1101101101;
    16'b0000000000001000: out_v[335] = 10'b0010101011;
    16'b0000000000100000: out_v[335] = 10'b0101101011;
    16'b0000001010100000: out_v[335] = 10'b0111110111;
    16'b0000000010100100: out_v[335] = 10'b1101001010;
    16'b0001001010100000: out_v[335] = 10'b1111101011;
    16'b0001000010100000: out_v[335] = 10'b0100100100;
    16'b0000100000000000: out_v[335] = 10'b1001100100;
    16'b0001000011100100: out_v[335] = 10'b0001101100;
    16'b0000000010100000: out_v[335] = 10'b0000011011;
    16'b0001000010100100: out_v[335] = 10'b0011000110;
    16'b0000000010101000: out_v[335] = 10'b1001011100;
    16'b0001000011101000: out_v[335] = 10'b0101001010;
    16'b0011100100101000: out_v[335] = 10'b1100010110;
    16'b0001000000100000: out_v[335] = 10'b0011101111;
    16'b0000100000100000: out_v[335] = 10'b1111000010;
    16'b0001001000100000: out_v[335] = 10'b1011011011;
    16'b0001000011100000: out_v[335] = 10'b1000011110;
    16'b0010100100101000: out_v[335] = 10'b0000100110;
    16'b0001100000100000: out_v[335] = 10'b1001100100;
    16'b0000000010001100: out_v[335] = 10'b1100100101;
    16'b0000100000101000: out_v[335] = 10'b0001110010;
    16'b0000101000100000: out_v[335] = 10'b0110000100;
    16'b0001000000001000: out_v[335] = 10'b1000001100;
    16'b0000000000101000: out_v[335] = 10'b0100100101;
    16'b0000001001100000: out_v[335] = 10'b1110101011;
    16'b0001001011100000: out_v[335] = 10'b0000011000;
    16'b0000001000100000: out_v[335] = 10'b0110110111;
    16'b0001000010101100: out_v[335] = 10'b1011011111;
    16'b0001100010100000: out_v[335] = 10'b1110100010;
    16'b0001000010101000: out_v[335] = 10'b0001010100;
    16'b0001001001100000: out_v[335] = 10'b1101110011;
    16'b0001000000101000: out_v[335] = 10'b1000000110;
    16'b0001000010001100: out_v[335] = 10'b1001110100;
    16'b0001101010100000: out_v[335] = 10'b0111010011;
    16'b0001101000100000: out_v[335] = 10'b1011100101;
    16'b0001100011100100: out_v[335] = 10'b1010011000;
    16'b0001100001100100: out_v[335] = 10'b0010001010;
    16'b0001100000100100: out_v[335] = 10'b1110101001;
    16'b0000000011100100: out_v[335] = 10'b0101010001;
    16'b0000100000100100: out_v[335] = 10'b0110100010;
    16'b0000100010100000: out_v[335] = 10'b1001010010;
    16'b0000000010101100: out_v[335] = 10'b1011011111;
    16'b0000100010000100: out_v[335] = 10'b1111101001;
    16'b0000000000100100: out_v[335] = 10'b1111110100;
    16'b0001000001100100: out_v[335] = 10'b0100011011;
    16'b0000100011100100: out_v[335] = 10'b1110100011;
    16'b0001100001100000: out_v[335] = 10'b1010110001;
    16'b0010100110001100: out_v[335] = 10'b0111101010;
    16'b0000100010000000: out_v[335] = 10'b1100010100;
    16'b0000100000001100: out_v[335] = 10'b0101111111;
    16'b0000100010001000: out_v[335] = 10'b0011010110;
    16'b0110100101101001: out_v[335] = 10'b1001010011;
    16'b0000100001000000: out_v[335] = 10'b1100101100;
    16'b0011100100100000: out_v[335] = 10'b0110010111;
    16'b0000100000001000: out_v[335] = 10'b0001111010;
    16'b0000100000000100: out_v[335] = 10'b0010111101;
    16'b0000100001100000: out_v[335] = 10'b0000011011;
    16'b0001100000000000: out_v[335] = 10'b1001110011;
    16'b0001100001100001: out_v[335] = 10'b1101010011;
    16'b0110000101101001: out_v[335] = 10'b1110111110;
    16'b0010100110001000: out_v[335] = 10'b0111011110;
    16'b0001100000000100: out_v[335] = 10'b0000110101;
    16'b0001100001000000: out_v[335] = 10'b0100111110;
    16'b0010100100001000: out_v[335] = 10'b1101011011;
    16'b0010000101101000: out_v[335] = 10'b1010101111;
    16'b0000100001101000: out_v[335] = 10'b0011111110;
    16'b0000100001001100: out_v[335] = 10'b0010101101;
    16'b0010100100001100: out_v[335] = 10'b1101101011;
    16'b0010100101101000: out_v[335] = 10'b0101010011;
    16'b0111100101100001: out_v[335] = 10'b1101011110;
    16'b0001100001000100: out_v[335] = 10'b1011110000;
    16'b0000100011001100: out_v[335] = 10'b1101011111;
    16'b0001100011100101: out_v[335] = 10'b1100011010;
    16'b0001100011000100: out_v[335] = 10'b0111010011;
    16'b0001100010000000: out_v[335] = 10'b1011101100;
    16'b0000100011000100: out_v[335] = 10'b1111010110;
    16'b0000000011000100: out_v[335] = 10'b1011110010;
    16'b0000100011100000: out_v[335] = 10'b0110010111;
    16'b0010000101110000: out_v[335] = 10'b1111011000;
    16'b0110000101110001: out_v[335] = 10'b0110101011;
    16'b0010100100110000: out_v[335] = 10'b0111111010;
    16'b0000100001110000: out_v[335] = 10'b1110010011;
    16'b0000100000110000: out_v[335] = 10'b0111100000;
    16'b0010000101110001: out_v[335] = 10'b0010111001;
    16'b0000100010110000: out_v[335] = 10'b1111111111;
    16'b0000000001100000: out_v[335] = 10'b1110000011;
    16'b0000000011001101: out_v[335] = 10'b0011111011;
    16'b0100000001101101: out_v[335] = 10'b1011111011;
    16'b0001000011001101: out_v[335] = 10'b0011111111;
    16'b0000000001100001: out_v[335] = 10'b0000101100;
    16'b0000000001100100: out_v[335] = 10'b1011010101;
    16'b0001000011000000: out_v[335] = 10'b0111001010;
    16'b0001000001000000: out_v[335] = 10'b1011110000;
    16'b0001000001000100: out_v[335] = 10'b1010010001;
    16'b0000000001101001: out_v[335] = 10'b0110001111;
    16'b0001000011001100: out_v[335] = 10'b1011010011;
    16'b0000000001000000: out_v[335] = 10'b1100011000;
    16'b0001000001000101: out_v[335] = 10'b0110011011;
    16'b0001000011000100: out_v[335] = 10'b0001011111;
    16'b0000000001001100: out_v[335] = 10'b1010000110;
    16'b0000000011001100: out_v[335] = 10'b1011001111;
    16'b0000000001000100: out_v[335] = 10'b0100110111;
    16'b0000000001001101: out_v[335] = 10'b0000101101;
    16'b0000000001101101: out_v[335] = 10'b0110101010;
    16'b0001000001001101: out_v[335] = 10'b0111110101;
    16'b0001000011001000: out_v[335] = 10'b0001110001;
    16'b0001000001001100: out_v[335] = 10'b0001001111;
    16'b0000000011001000: out_v[335] = 10'b1011000101;
    16'b0000000011001001: out_v[335] = 10'b0111010010;
    16'b0000000001000001: out_v[335] = 10'b0111001101;
    16'b0000000001000101: out_v[335] = 10'b1101101111;
    16'b0001000011001001: out_v[335] = 10'b0111100010;
    16'b0100000011001101: out_v[335] = 10'b0111100111;
    16'b0001100000001100: out_v[335] = 10'b1101001000;
    16'b0000000011101100: out_v[335] = 10'b1010100111;
    16'b0000100011101101: out_v[335] = 10'b0100111010;
    16'b0001100011101101: out_v[335] = 10'b0100111100;
    16'b0001100011001100: out_v[335] = 10'b1101110111;
    16'b0000100011101100: out_v[335] = 10'b1111000110;
    16'b0000000000001100: out_v[335] = 10'b0100101111;
    16'b0111000101100001: out_v[335] = 10'b1101000011;
    16'b0000100001000100: out_v[335] = 10'b1101011111;
    16'b0111000101101001: out_v[335] = 10'b1001001000;
    16'b0001100001001100: out_v[335] = 10'b1011100110;
    16'b0000100001100001: out_v[335] = 10'b1001010000;
    16'b0110100101100001: out_v[335] = 10'b1001010011;
    16'b0111100101101001: out_v[335] = 10'b1011001110;
    16'b0110000101100001: out_v[335] = 10'b1101000011;
    default: out_v[335] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010100011000000: out_v[336] = 10'b1011001101;
    16'b0000000011000000: out_v[336] = 10'b1110001101;
    16'b0000100001000000: out_v[336] = 10'b0100010110;
    16'b0000100011000000: out_v[336] = 10'b1100000101;
    16'b0000100000000000: out_v[336] = 10'b0011101101;
    16'b0000000000000000: out_v[336] = 10'b1011001110;
    16'b0010000011000000: out_v[336] = 10'b0100001001;
    16'b0000000010000000: out_v[336] = 10'b0000011011;
    16'b0010000010000000: out_v[336] = 10'b0101011011;
    16'b0000000001000000: out_v[336] = 10'b0000011001;
    16'b0000100010000000: out_v[336] = 10'b0101000101;
    16'b0010100010000000: out_v[336] = 10'b0111010100;
    16'b0010000000000000: out_v[336] = 10'b0010011010;
    16'b0010000001000000: out_v[336] = 10'b0100110010;
    16'b0010100000000000: out_v[336] = 10'b1101111001;
    16'b0010100001000000: out_v[336] = 10'b1010110011;
    16'b0000100111000000: out_v[336] = 10'b0101001011;
    16'b0010100111000000: out_v[336] = 10'b0010101101;
    16'b0000100110000000: out_v[336] = 10'b1101000000;
    16'b0000100101000000: out_v[336] = 10'b0111001010;
    16'b0000010000000000: out_v[336] = 10'b1000100010;
    16'b0000110000000000: out_v[336] = 10'b0101011000;
    16'b0010001000000000: out_v[336] = 10'b1011001110;
    16'b0010001001000000: out_v[336] = 10'b1011010011;
    16'b0010010011000000: out_v[336] = 10'b1000110111;
    16'b0000010001000000: out_v[336] = 10'b0110011100;
    16'b0000110001000000: out_v[336] = 10'b1010101000;
    16'b0000010011000000: out_v[336] = 10'b0110110000;
    16'b0010010001000000: out_v[336] = 10'b1001001110;
    16'b0000000110000000: out_v[336] = 10'b1111010000;
    16'b0000000111000000: out_v[336] = 10'b0001001010;
    16'b0000000101000000: out_v[336] = 10'b1011001011;
    16'b0010000000100000: out_v[336] = 10'b1111100011;
    16'b0000000000100000: out_v[336] = 10'b1110000110;
    16'b0000000000010000: out_v[336] = 10'b0011011010;
    16'b0000110011000000: out_v[336] = 10'b1100101011;
    default: out_v[336] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000100001000: out_v[337] = 10'b1100000001;
    16'b0001110000001110: out_v[337] = 10'b0111001110;
    16'b0000100100001000: out_v[337] = 10'b0010010111;
    16'b0000110100001101: out_v[337] = 10'b0000110111;
    16'b0011110000000110: out_v[337] = 10'b1110110110;
    16'b0010000000001110: out_v[337] = 10'b1000111001;
    16'b0010100000001110: out_v[337] = 10'b1100011111;
    16'b0000100100001001: out_v[337] = 10'b1011001100;
    16'b1001110100001100: out_v[337] = 10'b0110011110;
    16'b0001100000000110: out_v[337] = 10'b1110001001;
    16'b1000100100001111: out_v[337] = 10'b1010100111;
    16'b1001100000001110: out_v[337] = 10'b0010010101;
    16'b0001100100001110: out_v[337] = 10'b1011110011;
    16'b0001100000001000: out_v[337] = 10'b1000011011;
    16'b0001100000001110: out_v[337] = 10'b0011110000;
    16'b0000100100001101: out_v[337] = 10'b1110001010;
    16'b0011100000001110: out_v[337] = 10'b0111001110;
    16'b0011000000001110: out_v[337] = 10'b1111111001;
    16'b0001100100001100: out_v[337] = 10'b1010111001;
    16'b0000100000001110: out_v[337] = 10'b0111001011;
    16'b0000110000001110: out_v[337] = 10'b0011010110;
    16'b1000100100001100: out_v[337] = 10'b1100110111;
    16'b0000110000001111: out_v[337] = 10'b1110100011;
    16'b1000110100001101: out_v[337] = 10'b1100100111;
    16'b0001100000001010: out_v[337] = 10'b1010000011;
    16'b0011100000001111: out_v[337] = 10'b0111010010;
    16'b0001000000001110: out_v[337] = 10'b1101000011;
    16'b1000000100001001: out_v[337] = 10'b0000111111;
    16'b0000100000001111: out_v[337] = 10'b1010001001;
    16'b1001100100001110: out_v[337] = 10'b1010110111;
    16'b1000100100001101: out_v[337] = 10'b1110110001;
    16'b0000100000001100: out_v[337] = 10'b1101100011;
    16'b0001110000001111: out_v[337] = 10'b1110011010;
    16'b0001010000001110: out_v[337] = 10'b1111100111;
    16'b0000100100001100: out_v[337] = 10'b1011110111;
    16'b0000100000001010: out_v[337] = 10'b1101010001;
    16'b1000000100000001: out_v[337] = 10'b0001011011;
    16'b1000110100001111: out_v[337] = 10'b1001010111;
    16'b0011110000001110: out_v[337] = 10'b1110111101;
    16'b1001100100001111: out_v[337] = 10'b1111000111;
    16'b1011100000001110: out_v[337] = 10'b1011000111;
    16'b0001110100001110: out_v[337] = 10'b1110111010;
    16'b0001100100001000: out_v[337] = 10'b0001111011;
    16'b0001100000001100: out_v[337] = 10'b1111111011;
    16'b0001100000001111: out_v[337] = 10'b1011001011;
    16'b0000100000001000: out_v[337] = 10'b0111000011;
    16'b1001110100001111: out_v[337] = 10'b1010110011;
    16'b1000110100001100: out_v[337] = 10'b1011010100;
    16'b0001110000000110: out_v[337] = 10'b1111001111;
    16'b0000000000001110: out_v[337] = 10'b1011010011;
    16'b1000010000001000: out_v[337] = 10'b1111010101;
    16'b1000000000001000: out_v[337] = 10'b1111010001;
    16'b1000000000000000: out_v[337] = 10'b0100011011;
    16'b0000000000000000: out_v[337] = 10'b0001100111;
    16'b1000000000000001: out_v[337] = 10'b1100001001;
    16'b1000010000000000: out_v[337] = 10'b0110010110;
    16'b0000000000000001: out_v[337] = 10'b0010100100;
    16'b1000010100001000: out_v[337] = 10'b1001001110;
    16'b0000010000000000: out_v[337] = 10'b1001011011;
    16'b0000010000001000: out_v[337] = 10'b1001101110;
    16'b1000000100000000: out_v[337] = 10'b0011110000;
    16'b1000010100001001: out_v[337] = 10'b1010100101;
    16'b1000000100001000: out_v[337] = 10'b0101101010;
    16'b0000000000001000: out_v[337] = 10'b0011000100;
    16'b1000010100001100: out_v[337] = 10'b0011011110;
    16'b1000010100000000: out_v[337] = 10'b0000110100;
    16'b0100000000001000: out_v[337] = 10'b1100101111;
    16'b0001000000001101: out_v[337] = 10'b1011010110;
    16'b0000010000001101: out_v[337] = 10'b0001111110;
    16'b0000000000001101: out_v[337] = 10'b0010100110;
    16'b0001000000000000: out_v[337] = 10'b1000110010;
    16'b0000100000001101: out_v[337] = 10'b1100111110;
    16'b0000100100000101: out_v[337] = 10'b1010101111;
    16'b0000010000001001: out_v[337] = 10'b1010001111;
    16'b0001010000001101: out_v[337] = 10'b1001010110;
    16'b0000000100000001: out_v[337] = 10'b1101000001;
    16'b0000010000000101: out_v[337] = 10'b0110110101;
    16'b0001110100001101: out_v[337] = 10'b0000110110;
    16'b0001100100001101: out_v[337] = 10'b1001001110;
    16'b0000000000001100: out_v[337] = 10'b0011011111;
    16'b0000110000001101: out_v[337] = 10'b1010001001;
    16'b0001100100000101: out_v[337] = 10'b1111010110;
    16'b0000000000001001: out_v[337] = 10'b0010011010;
    16'b0001000000001001: out_v[337] = 10'b1011101010;
    16'b0001000000000101: out_v[337] = 10'b1010001110;
    16'b1001000100000000: out_v[337] = 10'b0110000100;
    16'b0001000000000001: out_v[337] = 10'b0010010111;
    16'b0000000000000101: out_v[337] = 10'b0001101110;
    16'b0000000100001101: out_v[337] = 10'b0111101010;
    16'b0001100000001101: out_v[337] = 10'b0110001100;
    16'b0000011000001101: out_v[337] = 10'b0101110110;
    16'b0000010000001100: out_v[337] = 10'b1001110111;
    16'b0000000000000100: out_v[337] = 10'b1000110110;
    16'b0001000100001101: out_v[337] = 10'b1011110110;
    16'b0000100100000001: out_v[337] = 10'b0010110100;
    16'b1001000100000001: out_v[337] = 10'b1111011100;
    16'b1001100100000101: out_v[337] = 10'b1111110000;
    16'b1001100100001101: out_v[337] = 10'b1000011110;
    16'b1001000100000101: out_v[337] = 10'b0011111011;
    16'b1001000000000000: out_v[337] = 10'b1110011100;
    16'b1001000100001100: out_v[337] = 10'b1111110001;
    16'b1000000100000101: out_v[337] = 10'b1001110011;
    16'b1001100100000000: out_v[337] = 10'b1001001110;
    16'b1001000100001000: out_v[337] = 10'b1001101010;
    16'b1000010100001101: out_v[337] = 10'b1100001011;
    16'b1000100100001000: out_v[337] = 10'b0111011110;
    16'b1001100100001000: out_v[337] = 10'b0011001010;
    16'b1001100100001010: out_v[337] = 10'b1011100110;
    16'b1000100100000001: out_v[337] = 10'b0010011111;
    16'b0000000100001001: out_v[337] = 10'b1001000011;
    16'b1001000000000100: out_v[337] = 10'b0010101010;
    16'b1001000100000100: out_v[337] = 10'b1110011101;
    16'b1000000000001001: out_v[337] = 10'b1101110001;
    16'b1000000100001101: out_v[337] = 10'b1110100010;
    16'b1001010100001100: out_v[337] = 10'b1111011110;
    16'b1000100100000000: out_v[337] = 10'b0010010101;
    16'b1000000000001100: out_v[337] = 10'b1100111000;
    16'b1000010000001101: out_v[337] = 10'b1111011000;
    16'b1000000000001101: out_v[337] = 10'b0101101010;
    16'b1001000000001100: out_v[337] = 10'b1111001010;
    16'b1000000100000100: out_v[337] = 10'b1011101100;
    16'b1001010100001000: out_v[337] = 10'b1111011110;
    16'b1001000000001000: out_v[337] = 10'b0110110110;
    16'b1000000100001100: out_v[337] = 10'b0001111110;
    16'b1001000100001001: out_v[337] = 10'b1100000011;
    16'b1000100100001001: out_v[337] = 10'b0010111110;
    16'b1001100100000010: out_v[337] = 10'b1100010100;
    16'b1000000000000100: out_v[337] = 10'b1001001011;
    16'b1000011100001001: out_v[337] = 10'b1100101001;
    16'b1000000000000101: out_v[337] = 10'b1100011010;
    16'b1001000100000010: out_v[337] = 10'b0111001010;
    16'b0000100000001011: out_v[337] = 10'b1101100110;
    16'b0000100000000011: out_v[337] = 10'b1101111010;
    16'b0000100100000011: out_v[337] = 10'b0000110011;
    16'b0000100100001010: out_v[337] = 10'b0011111011;
    16'b1000100100000011: out_v[337] = 10'b1011000111;
    16'b0001100000001011: out_v[337] = 10'b0010111110;
    16'b0000100100001011: out_v[337] = 10'b1101010011;
    16'b0000110000001001: out_v[337] = 10'b0101110100;
    16'b0000100000001001: out_v[337] = 10'b1001011011;
    16'b0000000100000011: out_v[337] = 10'b1101100001;
    16'b0100100100001011: out_v[337] = 10'b1110001101;
    16'b1000100100001011: out_v[337] = 10'b1000100110;
    16'b0000110000001011: out_v[337] = 10'b0001110011;
    16'b0100100100001001: out_v[337] = 10'b1011111111;
    16'b0000110100001011: out_v[337] = 10'b1111000011;
    16'b0001100100001011: out_v[337] = 10'b0100100011;
    16'b0100100000001011: out_v[337] = 10'b0011101100;
    16'b0100100100000011: out_v[337] = 10'b1011101110;
    16'b0000100000000001: out_v[337] = 10'b1101000011;
    16'b0010100100001011: out_v[337] = 10'b1100111100;
    16'b0000110100001001: out_v[337] = 10'b0011001100;
    16'b1000110100001011: out_v[337] = 10'b1000011110;
    16'b0000100100000010: out_v[337] = 10'b0110010010;
    16'b1100010100000001: out_v[337] = 10'b1011011101;
    16'b1001010000000100: out_v[337] = 10'b0110110011;
    16'b0000000100000000: out_v[337] = 10'b1011101001;
    16'b0000100100001111: out_v[337] = 10'b0101100010;
    16'b1100010000000101: out_v[337] = 10'b1110110111;
    16'b1000100100000010: out_v[337] = 10'b1101100010;
    16'b1000010100000001: out_v[337] = 10'b0111100101;
    16'b1100010100000101: out_v[337] = 10'b0010011111;
    16'b1100000100001101: out_v[337] = 10'b1010011110;
    16'b1001110100000010: out_v[337] = 10'b1100101100;
    16'b0000010100000001: out_v[337] = 10'b0010110011;
    16'b1000010000000001: out_v[337] = 10'b0010110001;
    16'b1001010100000000: out_v[337] = 10'b1010110101;
    16'b0001100000000000: out_v[337] = 10'b0111111011;
    16'b0001000100000001: out_v[337] = 10'b0011001010;
    16'b0001000100000000: out_v[337] = 10'b1110100011;
    16'b0001100100000001: out_v[337] = 10'b0011110010;
    16'b0011100000000111: out_v[337] = 10'b1110101011;
    16'b0011100000000010: out_v[337] = 10'b0011011000;
    16'b0001100100000000: out_v[337] = 10'b1110111111;
    16'b0001100000000011: out_v[337] = 10'b1100011001;
    16'b1001100100000001: out_v[337] = 10'b0001001101;
    16'b1000110100000101: out_v[337] = 10'b0111000010;
    16'b0011100000000011: out_v[337] = 10'b0111101110;
    16'b0000100000000000: out_v[337] = 10'b0010010001;
    16'b0001100000000111: out_v[337] = 10'b1010011011;
    16'b0000100000000010: out_v[337] = 10'b1011100011;
    16'b0001100000000001: out_v[337] = 10'b1101001001;
    16'b1000100100000101: out_v[337] = 10'b0111110001;
    16'b1001100100000100: out_v[337] = 10'b1101111110;
    16'b1000110100000001: out_v[337] = 10'b1001000011;
    16'b0001100000000010: out_v[337] = 10'b0110011111;
    16'b0000100000000101: out_v[337] = 10'b1011101100;
    16'b0000100000000111: out_v[337] = 10'b1101110010;
    16'b1001110100000100: out_v[337] = 10'b1101010101;
    16'b0000100100000000: out_v[337] = 10'b1000101100;
    16'b0000000000001011: out_v[337] = 10'b0010001100;
    16'b1000000000001011: out_v[337] = 10'b0111001100;
    16'b0000000000000011: out_v[337] = 10'b0010011100;
    16'b1000100000001011: out_v[337] = 10'b0001111110;
    16'b1000000000000011: out_v[337] = 10'b0100001111;
    16'b0000010100001000: out_v[337] = 10'b0100011011;
    16'b1000010000001001: out_v[337] = 10'b0111010100;
    16'b0000000100001011: out_v[337] = 10'b1101001011;
    16'b1000010100000100: out_v[337] = 10'b0111110000;
    16'b0000010100001101: out_v[337] = 10'b0110011011;
    16'b1000000100001011: out_v[337] = 10'b1000000111;
    16'b1000010100000101: out_v[337] = 10'b1000110001;
    16'b0000010100001001: out_v[337] = 10'b0011001100;
    16'b0000000100001100: out_v[337] = 10'b1110011100;
    16'b1000000100000011: out_v[337] = 10'b1000010110;
    default: out_v[337] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010000101000000: out_v[338] = 10'b1000001111;
    16'b0010100100000000: out_v[338] = 10'b0111010001;
    16'b0010100100000001: out_v[338] = 10'b0111000000;
    16'b0110100100000000: out_v[338] = 10'b0111011001;
    16'b0010100101000000: out_v[338] = 10'b1000001100;
    16'b0010000100000000: out_v[338] = 10'b0110110101;
    16'b0000100100000000: out_v[338] = 10'b1000100010;
    16'b0000100100010000: out_v[338] = 10'b0010100100;
    16'b0100100000000000: out_v[338] = 10'b0010110110;
    16'b0011100101000000: out_v[338] = 10'b0110010010;
    16'b0010000101010000: out_v[338] = 10'b0010000111;
    16'b0011100100000000: out_v[338] = 10'b1000011000;
    16'b0000100000000000: out_v[338] = 10'b1000100001;
    16'b0000100100000001: out_v[338] = 10'b1000100111;
    16'b0010100100010001: out_v[338] = 10'b0111001111;
    16'b0010000100010001: out_v[338] = 10'b0101010101;
    16'b0100100100000000: out_v[338] = 10'b1000001101;
    16'b0010000101010001: out_v[338] = 10'b0111000111;
    16'b0000100100010001: out_v[338] = 10'b0000100101;
    16'b0001100100000000: out_v[338] = 10'b1000100001;
    16'b0000100101000000: out_v[338] = 10'b1011011001;
    16'b0010000001000000: out_v[338] = 10'b1100011110;
    16'b0111100100000000: out_v[338] = 10'b0000011110;
    16'b0010000000000000: out_v[338] = 10'b1010010101;
    16'b0010100000000000: out_v[338] = 10'b0010011101;
    16'b0010000100010000: out_v[338] = 10'b1010101110;
    16'b0011000101000000: out_v[338] = 10'b1101000100;
    16'b0010100101010001: out_v[338] = 10'b1111010011;
    16'b0000000100000000: out_v[338] = 10'b1001100000;
    16'b0110100000000000: out_v[338] = 10'b1011000101;
    16'b0011000100000000: out_v[338] = 10'b1001100110;
    16'b0011100001000000: out_v[338] = 10'b0110110111;
    16'b0011100000000000: out_v[338] = 10'b1001011111;
    16'b0001000100000000: out_v[338] = 10'b0000111010;
    16'b0001000000000000: out_v[338] = 10'b1001011110;
    16'b0001100001000000: out_v[338] = 10'b0001010011;
    16'b0001100000000000: out_v[338] = 10'b0010110001;
    16'b0001000001000000: out_v[338] = 10'b0000000100;
    16'b0001000101000000: out_v[338] = 10'b1111010001;
    16'b0000000000000000: out_v[338] = 10'b0001110010;
    16'b0001000100010000: out_v[338] = 10'b0010001000;
    16'b0001000101010000: out_v[338] = 10'b0111011100;
    16'b0001000100010001: out_v[338] = 10'b1001000101;
    16'b0011000101010000: out_v[338] = 10'b1101000100;
    16'b0111100001000000: out_v[338] = 10'b0110011110;
    16'b0010100001000000: out_v[338] = 10'b1100001111;
    16'b0000000001000000: out_v[338] = 10'b1101001010;
    16'b0010000000010001: out_v[338] = 10'b1101000111;
    16'b0100100001000000: out_v[338] = 10'b0011001011;
    16'b0010100000010000: out_v[338] = 10'b1010100011;
    16'b0110100001000000: out_v[338] = 10'b0110100110;
    16'b0001000101010001: out_v[338] = 10'b1011110001;
    16'b0010000000010000: out_v[338] = 10'b0011001010;
    16'b0011000001010000: out_v[338] = 10'b1010010011;
    16'b0011000101010001: out_v[338] = 10'b0110010001;
    16'b0010000001010000: out_v[338] = 10'b0101111110;
    16'b0010000001010001: out_v[338] = 10'b0101111110;
    16'b0011100101010000: out_v[338] = 10'b1110000101;
    16'b0010100101010000: out_v[338] = 10'b1000011100;
    16'b0011000001000000: out_v[338] = 10'b0101101011;
    16'b0001000001010001: out_v[338] = 10'b0100011111;
    16'b0001000000010001: out_v[338] = 10'b1110001110;
    16'b0001000001000001: out_v[338] = 10'b1100101011;
    16'b0001000000010000: out_v[338] = 10'b0010111011;
    16'b0011100101010001: out_v[338] = 10'b0101001110;
    16'b0001000001010000: out_v[338] = 10'b1100010011;
    16'b0011000001010001: out_v[338] = 10'b1001101000;
    16'b0010100001010000: out_v[338] = 10'b1110010101;
    16'b0001000100000001: out_v[338] = 10'b0101011011;
    16'b0000000100010000: out_v[338] = 10'b0010111000;
    16'b0011100100010001: out_v[338] = 10'b1100011010;
    16'b0011000100010000: out_v[338] = 10'b0010111010;
    16'b0111100100010000: out_v[338] = 10'b1111111010;
    16'b0011100100010000: out_v[338] = 10'b1011011011;
    16'b0011000100010001: out_v[338] = 10'b1110100010;
    16'b0111100000000000: out_v[338] = 10'b0000011000;
    16'b0001100100010000: out_v[338] = 10'b0101100011;
    16'b0011100100000001: out_v[338] = 10'b0011001010;
    16'b0000000100010001: out_v[338] = 10'b0101011111;
    16'b0001100100010001: out_v[338] = 10'b1010110111;
    16'b0011000100000001: out_v[338] = 10'b1010110010;
    16'b0101100100000000: out_v[338] = 10'b1111110011;
    16'b0111100100010001: out_v[338] = 10'b1010100101;
    16'b0001000000000001: out_v[338] = 10'b0010010001;
    16'b0011000000000000: out_v[338] = 10'b1001100010;
    16'b0010100000010001: out_v[338] = 10'b1110000101;
    16'b0000000000000001: out_v[338] = 10'b0011011110;
    16'b0011000000000001: out_v[338] = 10'b1011100000;
    16'b0010100001000001: out_v[338] = 10'b0010111010;
    16'b0010000000000001: out_v[338] = 10'b1010011100;
    16'b0010100000000001: out_v[338] = 10'b0011000110;
    16'b0010100001010001: out_v[338] = 10'b0110010110;
    16'b0000000000010000: out_v[338] = 10'b1011011010;
    16'b0011000000010001: out_v[338] = 10'b0001110011;
    16'b0011100000000001: out_v[338] = 10'b1001111100;
    16'b0010100100010000: out_v[338] = 10'b1101110110;
    16'b0000100001000000: out_v[338] = 10'b1100101010;
    16'b0001100101000000: out_v[338] = 10'b0110000001;
    16'b0001100100000001: out_v[338] = 10'b1100101111;
    16'b0101100000000000: out_v[338] = 10'b1111110111;
    16'b0000000101000000: out_v[338] = 10'b1101001110;
    16'b0000000001010001: out_v[338] = 10'b1010011110;
    16'b0000000001010000: out_v[338] = 10'b1110000110;
    16'b0010000100000001: out_v[338] = 10'b0101011110;
    16'b0001000101000001: out_v[338] = 10'b0110000011;
    16'b0000000100000001: out_v[338] = 10'b1010101010;
    16'b0011100101000001: out_v[338] = 10'b1011010111;
    16'b0011000101000001: out_v[338] = 10'b1001100110;
    default: out_v[338] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100000000000010: out_v[339] = 10'b0110010101;
    16'b0010000000000010: out_v[339] = 10'b0100001011;
    16'b1010100000000010: out_v[339] = 10'b1000111111;
    16'b1010000001000000: out_v[339] = 10'b0111001011;
    16'b0010000001000000: out_v[339] = 10'b0000110100;
    16'b0100000000000000: out_v[339] = 10'b0000110101;
    16'b1010000000000000: out_v[339] = 10'b1111001000;
    16'b1100000000000000: out_v[339] = 10'b1000110111;
    16'b1010100000000000: out_v[339] = 10'b1011000111;
    16'b0010000000000000: out_v[339] = 10'b0111001110;
    16'b0110000000000000: out_v[339] = 10'b0001101110;
    16'b0010000001000010: out_v[339] = 10'b1001001111;
    16'b0110000001000010: out_v[339] = 10'b0100001010;
    16'b0110000001000000: out_v[339] = 10'b0100010000;
    16'b1110000000000000: out_v[339] = 10'b1011010000;
    16'b0000000001000000: out_v[339] = 10'b1000100110;
    16'b1010000001000010: out_v[339] = 10'b1001011101;
    16'b0000000000000000: out_v[339] = 10'b1001001010;
    16'b1010100001000000: out_v[339] = 10'b1001111101;
    16'b1000000001000000: out_v[339] = 10'b1110011001;
    16'b1000000001000010: out_v[339] = 10'b0111011011;
    16'b0010100000000000: out_v[339] = 10'b1101000111;
    16'b0100000001000000: out_v[339] = 10'b0110011010;
    16'b1010100001000010: out_v[339] = 10'b0101010011;
    16'b0000000000000010: out_v[339] = 10'b0100001110;
    16'b1000000000000000: out_v[339] = 10'b1100011001;
    16'b1010000000000010: out_v[339] = 10'b1110110110;
    16'b0000100000000000: out_v[339] = 10'b1101100000;
    16'b0110000000000010: out_v[339] = 10'b0010101000;
    16'b1110000001000000: out_v[339] = 10'b1100001011;
    16'b1110000001000010: out_v[339] = 10'b0101100001;
    16'b0100000001000010: out_v[339] = 10'b1101010101;
    16'b0010100000000010: out_v[339] = 10'b0111001011;
    16'b0000000001000010: out_v[339] = 10'b0100101100;
    16'b0100000000100010: out_v[339] = 10'b1111000010;
    16'b0110000000100010: out_v[339] = 10'b0011101001;
    16'b0000000000100010: out_v[339] = 10'b0000111000;
    16'b1100000000100010: out_v[339] = 10'b1111000010;
    16'b1100000000000010: out_v[339] = 10'b1010111100;
    16'b1100000001000010: out_v[339] = 10'b0110010100;
    16'b0100000000100000: out_v[339] = 10'b0011010000;
    16'b1100000001000000: out_v[339] = 10'b0011101010;
    16'b0000110000000000: out_v[339] = 10'b0011111110;
    16'b0000010000000000: out_v[339] = 10'b1000101111;
    16'b1110000000000010: out_v[339] = 10'b1001110011;
    16'b0000000100000000: out_v[339] = 10'b0111001010;
    16'b0110000100000000: out_v[339] = 10'b0100010101;
    16'b0010000100000000: out_v[339] = 10'b1001101010;
    16'b0100000100000000: out_v[339] = 10'b1011010101;
    16'b0000000000100000: out_v[339] = 10'b0011110001;
    16'b0100000010100010: out_v[339] = 10'b1000111100;
    16'b0100000010000000: out_v[339] = 10'b1111100011;
    16'b0100000010100000: out_v[339] = 10'b0100101111;
    16'b0100110000000000: out_v[339] = 10'b0110001010;
    16'b0100100000000000: out_v[339] = 10'b0111000010;
    16'b0100100000000010: out_v[339] = 10'b0010111100;
    16'b0100100001000010: out_v[339] = 10'b0101001010;
    default: out_v[339] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010001000000000: out_v[340] = 10'b0011110100;
    16'b0000001000000100: out_v[340] = 10'b0010001110;
    16'b0100101000000100: out_v[340] = 10'b1101000111;
    16'b0100000000000000: out_v[340] = 10'b1001011000;
    16'b0000001000000000: out_v[340] = 10'b0011010110;
    16'b0100000000000100: out_v[340] = 10'b1011010011;
    16'b0100001000000100: out_v[340] = 10'b0010010001;
    16'b0000000000000010: out_v[340] = 10'b1001000110;
    16'b0000001010000100: out_v[340] = 10'b1101011001;
    16'b0100001000000000: out_v[340] = 10'b1010100111;
    16'b0010001000000100: out_v[340] = 10'b0111000111;
    16'b0010000000000100: out_v[340] = 10'b1111010010;
    16'b0100000000000110: out_v[340] = 10'b1000000011;
    16'b0100000000000010: out_v[340] = 10'b0001100001;
    16'b0110000000000100: out_v[340] = 10'b1100000101;
    16'b0000001000000110: out_v[340] = 10'b1101011000;
    16'b0000101010000100: out_v[340] = 10'b1000110111;
    16'b0000101000000100: out_v[340] = 10'b0010100100;
    16'b0000001010000000: out_v[340] = 10'b1001110000;
    16'b0000000000000110: out_v[340] = 10'b0010000101;
    16'b0100100000000000: out_v[340] = 10'b0010110011;
    16'b0100001000000110: out_v[340] = 10'b0110111111;
    16'b0100101000000000: out_v[340] = 10'b1111011001;
    16'b0110001000000100: out_v[340] = 10'b0111111000;
    16'b0110000000000000: out_v[340] = 10'b1001001001;
    16'b0010000000000000: out_v[340] = 10'b0010101110;
    16'b0000000000000100: out_v[340] = 10'b1010001110;
    16'b0000000000000000: out_v[340] = 10'b0010100111;
    16'b0110000000000110: out_v[340] = 10'b1101010111;
    16'b0100101010000100: out_v[340] = 10'b0010101111;
    16'b0000001010000110: out_v[340] = 10'b0100011010;
    16'b0100001010000100: out_v[340] = 10'b1100001001;
    16'b0010001010000100: out_v[340] = 10'b1100010101;
    16'b0000000010000100: out_v[340] = 10'b0000001110;
    16'b0000000010000000: out_v[340] = 10'b1100101100;
    16'b0010000010000100: out_v[340] = 10'b0001011110;
    16'b0000001010000010: out_v[340] = 10'b0100100011;
    16'b0000001000000010: out_v[340] = 10'b0000101010;
    16'b0010000010000000: out_v[340] = 10'b1100000010;
    16'b1000000010000110: out_v[340] = 10'b1001100110;
    16'b0000000010000010: out_v[340] = 10'b0110101001;
    16'b0000000010000110: out_v[340] = 10'b0011011100;
    16'b0100000010000100: out_v[340] = 10'b1101010100;
    16'b0100000010000110: out_v[340] = 10'b1101001010;
    16'b0100000010000000: out_v[340] = 10'b1011100110;
    16'b0100000010000010: out_v[340] = 10'b1111100110;
    16'b1000000000000110: out_v[340] = 10'b0001010101;
    16'b0000000010100000: out_v[340] = 10'b1111001100;
    16'b0010000000000110: out_v[340] = 10'b0110111101;
    16'b0000000000100000: out_v[340] = 10'b0010110000;
    16'b1000000000000010: out_v[340] = 10'b0000101100;
    16'b0010001000000010: out_v[340] = 10'b1010001011;
    16'b0010001010000110: out_v[340] = 10'b0111100101;
    16'b0010000010000010: out_v[340] = 10'b1110100000;
    16'b0010001000000110: out_v[340] = 10'b0001101001;
    16'b0010000010000110: out_v[340] = 10'b0011100001;
    16'b0010001010000010: out_v[340] = 10'b0001100111;
    16'b0010001010000000: out_v[340] = 10'b0010110011;
    16'b0100001010000110: out_v[340] = 10'b1011001100;
    16'b0110000010000000: out_v[340] = 10'b1111100010;
    16'b0110000010000100: out_v[340] = 10'b0001111110;
    16'b0110001010000000: out_v[340] = 10'b0000111101;
    16'b0100101010000000: out_v[340] = 10'b0000011001;
    16'b0100001010000000: out_v[340] = 10'b0010110110;
    16'b0100100010000000: out_v[340] = 10'b1011001110;
    16'b0110001010000100: out_v[340] = 10'b1001011111;
    16'b0010101010000100: out_v[340] = 10'b1101110110;
    16'b0000100010000100: out_v[340] = 10'b1101100000;
    16'b0000101010000000: out_v[340] = 10'b1110011010;
    16'b0010100010000100: out_v[340] = 10'b0100011001;
    16'b0100100010000100: out_v[340] = 10'b0011100110;
    16'b0000001010100000: out_v[340] = 10'b1011001100;
    16'b0000001000100000: out_v[340] = 10'b0001110011;
    16'b0000001010100100: out_v[340] = 10'b1100011011;
    16'b0000001110100100: out_v[340] = 10'b1101010011;
    16'b0110101000000100: out_v[340] = 10'b1000100111;
    16'b0000100000000100: out_v[340] = 10'b0111100010;
    16'b0010101010000000: out_v[340] = 10'b1000001101;
    16'b0000100010000000: out_v[340] = 10'b1111011110;
    16'b0010100010000000: out_v[340] = 10'b0111001011;
    16'b0100000000001100: out_v[340] = 10'b1101101111;
    16'b0100000010001100: out_v[340] = 10'b1101001011;
    default: out_v[340] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000100000000100: out_v[341] = 10'b1001001010;
    16'b0000100000000101: out_v[341] = 10'b0110001111;
    16'b0000100000001001: out_v[341] = 10'b0000000101;
    16'b0000000000000100: out_v[341] = 10'b0001010100;
    16'b0000100000001000: out_v[341] = 10'b1000111101;
    16'b0000100000000001: out_v[341] = 10'b0011101101;
    16'b0000100000000000: out_v[341] = 10'b0110100010;
    16'b0000000000001000: out_v[341] = 10'b0011011110;
    16'b0000100000001101: out_v[341] = 10'b0110100110;
    16'b0000000000001001: out_v[341] = 10'b0000101111;
    16'b0000000000000000: out_v[341] = 10'b1100110010;
    16'b0000100000001100: out_v[341] = 10'b1100100101;
    16'b0000000000000101: out_v[341] = 10'b1101010110;
    16'b0000000000001100: out_v[341] = 10'b1101010000;
    16'b0000000000000001: out_v[341] = 10'b1010011110;
    16'b0000000000001101: out_v[341] = 10'b0100100000;
    16'b0000110000000000: out_v[341] = 10'b1010010100;
    16'b0000010000000000: out_v[341] = 10'b1011100000;
    default: out_v[341] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000100011000: out_v[342] = 10'b0010100101;
    16'b0000000000011001: out_v[342] = 10'b1000101011;
    16'b0000000101010001: out_v[342] = 10'b1010100011;
    16'b0000000100010000: out_v[342] = 10'b0101110010;
    16'b0000000000011000: out_v[342] = 10'b1001111011;
    16'b0100001101011000: out_v[342] = 10'b0000011011;
    16'b0000000100011001: out_v[342] = 10'b1010101110;
    16'b0000000101000001: out_v[342] = 10'b1010110111;
    16'b0100001101000001: out_v[342] = 10'b0011101110;
    16'b0000000001011001: out_v[342] = 10'b1011000111;
    16'b0100000101011001: out_v[342] = 10'b1011000111;
    16'b0000000101011001: out_v[342] = 10'b0100111111;
    16'b0000000101000000: out_v[342] = 10'b0011001001;
    16'b0000000101010000: out_v[342] = 10'b1110110000;
    16'b0000000100010001: out_v[342] = 10'b1110011000;
    16'b0000000101011000: out_v[342] = 10'b1111100010;
    16'b0000000100000001: out_v[342] = 10'b0111101010;
    16'b0100001101011001: out_v[342] = 10'b0000100001;
    16'b0100001101000000: out_v[342] = 10'b0001111100;
    16'b0000000001011000: out_v[342] = 10'b1001011000;
    16'b0100001101010001: out_v[342] = 10'b1101110110;
    16'b0100001101100001: out_v[342] = 10'b1001101100;
    16'b0100001101111001: out_v[342] = 10'b1110111011;
    16'b0000000100000000: out_v[342] = 10'b0001001111;
    16'b0100001101100101: out_v[342] = 10'b1100110001;
    16'b0100000101010001: out_v[342] = 10'b1001111110;
    16'b0000000000010000: out_v[342] = 10'b1100011001;
    16'b0100000101000001: out_v[342] = 10'b1111111010;
    16'b0100000101000000: out_v[342] = 10'b1010111101;
    16'b0100001001100101: out_v[342] = 10'b0011011001;
    16'b0100001101111101: out_v[342] = 10'b1011100010;
    16'b0000000000000000: out_v[342] = 10'b0010001110;
    16'b0000000000001000: out_v[342] = 10'b1100110010;
    16'b0000000001001000: out_v[342] = 10'b1100110000;
    16'b0100000000000000: out_v[342] = 10'b1100100111;
    16'b0100001001000000: out_v[342] = 10'b1101000100;
    16'b0000000001000000: out_v[342] = 10'b1000100101;
    16'b0100001100000000: out_v[342] = 10'b0111110000;
    16'b0000000000000001: out_v[342] = 10'b0010101100;
    16'b0000000001000001: out_v[342] = 10'b0111010110;
    16'b0100001000000000: out_v[342] = 10'b0001000111;
    16'b0000000011000000: out_v[342] = 10'b1010110011;
    16'b0000000010000000: out_v[342] = 10'b1011101110;
    16'b0000000001000010: out_v[342] = 10'b1010000010;
    16'b0100000001000000: out_v[342] = 10'b0101000110;
    16'b0000000001100100: out_v[342] = 10'b1100010010;
    16'b0100001001011000: out_v[342] = 10'b1010001010;
    16'b0000000101001000: out_v[342] = 10'b0100100111;
    16'b0000000001000100: out_v[342] = 10'b0101111111;
    16'b0000000001010000: out_v[342] = 10'b0111001010;
    16'b0000000101100100: out_v[342] = 10'b1000001101;
    16'b0000000100001000: out_v[342] = 10'b1110000000;
    16'b0000000101000100: out_v[342] = 10'b0001001000;
    16'b0100001100010000: out_v[342] = 10'b0110011011;
    16'b0000000000100100: out_v[342] = 10'b1001010011;
    16'b0000000100100000: out_v[342] = 10'b0001111101;
    16'b0000000000100000: out_v[342] = 10'b1111110111;
    16'b0000010000011000: out_v[342] = 10'b0001111110;
    16'b0000010100011000: out_v[342] = 10'b1001101100;
    16'b0000010000010000: out_v[342] = 10'b0010100100;
    16'b0000010100000000: out_v[342] = 10'b1100010100;
    16'b0000010000001000: out_v[342] = 10'b1110010001;
    16'b0000010101010000: out_v[342] = 10'b1000100011;
    16'b0000010100010000: out_v[342] = 10'b0011010001;
    16'b0000000111011000: out_v[342] = 10'b1010111111;
    16'b0000000001011010: out_v[342] = 10'b1111100011;
    16'b0000000100011010: out_v[342] = 10'b1000111110;
    16'b0100001101010000: out_v[342] = 10'b0111010011;
    16'b0000000010001000: out_v[342] = 10'b1001110001;
    16'b0000000010011000: out_v[342] = 10'b1010010010;
    16'b0100001101000010: out_v[342] = 10'b1111110100;
    16'b0000000011011000: out_v[342] = 10'b0111000010;
    16'b0100001101010010: out_v[342] = 10'b1110100000;
    16'b0000000101000010: out_v[342] = 10'b0011111001;
    16'b0000000000011010: out_v[342] = 10'b0111101011;
    16'b0000000100010010: out_v[342] = 10'b1011111111;
    16'b0000000111010000: out_v[342] = 10'b0100111001;
    16'b0000000101010010: out_v[342] = 10'b0110101101;
    16'b0000000101011010: out_v[342] = 10'b1000110111;
    16'b0100000101010000: out_v[342] = 10'b0111110101;
    16'b0000000000010010: out_v[342] = 10'b1101011011;
    16'b0000000000001010: out_v[342] = 10'b0111100010;
    16'b0000000100111101: out_v[342] = 10'b1111111011;
    16'b0000000101111100: out_v[342] = 10'b1110001110;
    16'b0000000100011100: out_v[342] = 10'b0001101111;
    16'b0000000100000100: out_v[342] = 10'b1011010110;
    16'b0000000100100100: out_v[342] = 10'b0010001111;
    16'b0000000100111000: out_v[342] = 10'b0110010011;
    16'b0000000000111100: out_v[342] = 10'b1110000100;
    16'b0000000100111100: out_v[342] = 10'b0111101100;
    16'b0001000100111100: out_v[342] = 10'b0001010000;
    16'b0000000100101100: out_v[342] = 10'b1011101110;
    16'b0000000100001100: out_v[342] = 10'b1100100101;
    16'b0000000000001001: out_v[342] = 10'b0110000000;
    default: out_v[342] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000100000001000: out_v[343] = 10'b1010110010;
    16'b0000100100000010: out_v[343] = 10'b0101011001;
    16'b0010110100000010: out_v[343] = 10'b1101101010;
    16'b0000100101001010: out_v[343] = 10'b0100010001;
    16'b0000110100001010: out_v[343] = 10'b1010110001;
    16'b0000100000000010: out_v[343] = 10'b0000101111;
    16'b0000110100000010: out_v[343] = 10'b0101100000;
    16'b0010110100000000: out_v[343] = 10'b0001011011;
    16'b0000010100000010: out_v[343] = 10'b1001110100;
    16'b0000100100001010: out_v[343] = 10'b0010001101;
    16'b0000100100000000: out_v[343] = 10'b0111110000;
    16'b0000100100001000: out_v[343] = 10'b0011100011;
    16'b0000100000000000: out_v[343] = 10'b0100110010;
    16'b0010110100001010: out_v[343] = 10'b1010010001;
    16'b0010011100000010: out_v[343] = 10'b0011110101;
    16'b0010010000000010: out_v[343] = 10'b0011100100;
    16'b0000000100000010: out_v[343] = 10'b1100110011;
    16'b0000000000000010: out_v[343] = 10'b0001010101;
    16'b0010010000000000: out_v[343] = 10'b0010011111;
    16'b0010011100000000: out_v[343] = 10'b1100011011;
    16'b0010010100000000: out_v[343] = 10'b0000110111;
    16'b0000010000000010: out_v[343] = 10'b1100100001;
    16'b0010010100000010: out_v[343] = 10'b1010010010;
    16'b0000100000001010: out_v[343] = 10'b0110011000;
    16'b0000000100001000: out_v[343] = 10'b0110010011;
    16'b0000110000000010: out_v[343] = 10'b1010110001;
    16'b0000000000000000: out_v[343] = 10'b1000000010;
    16'b0000000100000000: out_v[343] = 10'b1000100110;
    16'b0000000101000000: out_v[343] = 10'b0110111000;
    16'b0000000000001000: out_v[343] = 10'b0011110000;
    16'b0000100100010000: out_v[343] = 10'b0000001110;
    16'b0000100001000000: out_v[343] = 10'b1011001101;
    16'b0000100001001000: out_v[343] = 10'b0010101001;
    16'b0000100101001000: out_v[343] = 10'b1001001010;
    16'b0000100000011000: out_v[343] = 10'b1000001101;
    16'b0000000101001000: out_v[343] = 10'b0011101100;
    16'b0000000100010000: out_v[343] = 10'b0010010100;
    16'b0000100101000000: out_v[343] = 10'b1100000010;
    16'b0000101010000000: out_v[343] = 10'b1100100101;
    16'b0000101000000000: out_v[343] = 10'b1110100101;
    16'b0000110100001000: out_v[343] = 10'b0110001110;
    16'b0000100100011000: out_v[343] = 10'b0011000100;
    16'b0000101100001000: out_v[343] = 10'b0011101000;
    16'b0000000100011000: out_v[343] = 10'b1011101110;
    16'b0000000001000000: out_v[343] = 10'b0010001100;
    16'b0000100000010000: out_v[343] = 10'b1011000111;
    16'b0000101110000000: out_v[343] = 10'b1010001110;
    16'b0000101100000000: out_v[343] = 10'b0100110001;
    16'b0000000001001000: out_v[343] = 10'b0001110011;
    16'b0000000000001010: out_v[343] = 10'b0010011100;
    16'b0100000100001000: out_v[343] = 10'b1110101010;
    16'b0100100100001000: out_v[343] = 10'b0100111100;
    16'b0000000100001010: out_v[343] = 10'b0001010101;
    16'b0000110000001000: out_v[343] = 10'b0000111001;
    16'b0100000000001000: out_v[343] = 10'b1001011101;
    16'b0000110000001010: out_v[343] = 10'b1011010010;
    16'b0000010100001010: out_v[343] = 10'b1100110000;
    16'b0000010000001010: out_v[343] = 10'b1100001010;
    16'b0010110000001010: out_v[343] = 10'b0001010101;
    16'b0010010100001010: out_v[343] = 10'b1100010011;
    16'b0110110000001010: out_v[343] = 10'b0011111011;
    16'b0010110000001000: out_v[343] = 10'b1001100110;
    16'b0000100101000010: out_v[343] = 10'b1001011101;
    16'b0000110101001010: out_v[343] = 10'b0001011000;
    16'b0000111110001010: out_v[343] = 10'b0111100010;
    16'b0000000101001010: out_v[343] = 10'b1011001110;
    16'b0000100001001010: out_v[343] = 10'b0111001111;
    16'b0000010101001010: out_v[343] = 10'b0111011110;
    16'b1010010100001000: out_v[343] = 10'b0001111010;
    16'b1000010100001000: out_v[343] = 10'b0111110001;
    16'b0100100000001000: out_v[343] = 10'b0010100110;
    16'b1000000100001000: out_v[343] = 10'b1110000111;
    16'b1000000100001010: out_v[343] = 10'b0010001110;
    16'b0100010100001000: out_v[343] = 10'b0101011011;
    16'b0000010100001000: out_v[343] = 10'b0111100011;
    16'b0110110100001000: out_v[343] = 10'b0011001010;
    16'b1000010100001010: out_v[343] = 10'b1000000011;
    16'b0100110000001000: out_v[343] = 10'b1111101100;
    16'b0100110100001000: out_v[343] = 10'b0011101011;
    16'b1000000100000000: out_v[343] = 10'b1101100110;
    16'b0010010100001000: out_v[343] = 10'b1100011100;
    16'b0000010000001000: out_v[343] = 10'b0111001101;
    16'b0000010100000000: out_v[343] = 10'b0011010101;
    16'b0010110100001000: out_v[343] = 10'b1011011011;
    16'b0110110000001000: out_v[343] = 10'b0110101010;
    16'b0000110000000000: out_v[343] = 10'b0101001100;
    16'b0000110100000000: out_v[343] = 10'b0110011011;
    default: out_v[343] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000010000000: out_v[344] = 10'b1001100010;
    16'b0100000011000000: out_v[344] = 10'b1100000101;
    16'b0100000111000000: out_v[344] = 10'b0110110000;
    16'b0100000111000010: out_v[344] = 10'b1000010011;
    16'b0100000000000000: out_v[344] = 10'b0101011010;
    16'b0100000110000010: out_v[344] = 10'b0001101001;
    16'b0100000010000010: out_v[344] = 10'b1000000111;
    16'b0000000110000000: out_v[344] = 10'b0101011101;
    16'b0000000100000000: out_v[344] = 10'b1000001111;
    16'b0100000110000000: out_v[344] = 10'b0101101001;
    16'b0000000011000000: out_v[344] = 10'b1011001100;
    16'b0100000010000000: out_v[344] = 10'b1010000111;
    16'b0100000001000000: out_v[344] = 10'b0010011101;
    16'b0000000110000010: out_v[344] = 10'b1101110011;
    16'b0001000010000000: out_v[344] = 10'b0100011111;
    16'b0100000100000010: out_v[344] = 10'b0110010001;
    16'b0000000111000010: out_v[344] = 10'b0001100101;
    16'b0000000111000000: out_v[344] = 10'b0010001011;
    16'b0100000100000000: out_v[344] = 10'b1011100010;
    16'b0100000101000000: out_v[344] = 10'b0110011111;
    16'b0101000010000000: out_v[344] = 10'b0010110111;
    16'b0000000000000000: out_v[344] = 10'b0111110010;
    16'b0100000011000010: out_v[344] = 10'b1100000011;
    16'b0000000001000000: out_v[344] = 10'b0100110010;
    16'b0001000000000000: out_v[344] = 10'b0001000000;
    16'b0101000000000000: out_v[344] = 10'b0001100000;
    16'b0000000010000100: out_v[344] = 10'b1110000010;
    16'b0001000110000000: out_v[344] = 10'b1101000100;
    16'b0000100010000000: out_v[344] = 10'b0010111110;
    16'b0000000011000100: out_v[344] = 10'b1100001010;
    16'b0000000000000100: out_v[344] = 10'b0000001111;
    16'b0000000111000100: out_v[344] = 10'b1101011111;
    16'b0000000010000001: out_v[344] = 10'b1000100000;
    16'b0000000010000010: out_v[344] = 10'b0100111100;
    16'b0000000000000001: out_v[344] = 10'b1110010000;
    16'b0000000000000010: out_v[344] = 10'b0100011100;
    16'b0100000000000010: out_v[344] = 10'b0111010010;
    16'b0000000101000000: out_v[344] = 10'b1100011101;
    16'b0000000100000010: out_v[344] = 10'b0011000110;
    16'b0000000011000010: out_v[344] = 10'b0010111110;
    16'b0101000100000000: out_v[344] = 10'b0001101100;
    16'b0001000100000000: out_v[344] = 10'b1001110100;
    16'b0101000110000000: out_v[344] = 10'b1011011111;
    16'b0000000010000101: out_v[344] = 10'b0110011011;
    16'b0000000000010001: out_v[344] = 10'b1111010111;
    16'b0100000011000100: out_v[344] = 10'b0110100000;
    16'b0100000000000100: out_v[344] = 10'b0000010110;
    16'b0000000000000101: out_v[344] = 10'b1011001110;
    16'b0100000000010000: out_v[344] = 10'b1101101110;
    16'b0100000000010010: out_v[344] = 10'b1110001011;
    16'b0100000010000001: out_v[344] = 10'b0110001111;
    16'b0000000010000011: out_v[344] = 10'b0100111001;
    16'b0100000010000011: out_v[344] = 10'b1101100100;
    default: out_v[344] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010000001000011: out_v[345] = 10'b1000011111;
    16'b0000000101000010: out_v[345] = 10'b0011100110;
    16'b0110010101100010: out_v[345] = 10'b0000010111;
    16'b0110010101100011: out_v[345] = 10'b0001001111;
    16'b0110000001000011: out_v[345] = 10'b0000001011;
    16'b0000010100100010: out_v[345] = 10'b1010100100;
    16'b0110000101100010: out_v[345] = 10'b0111111001;
    16'b0010000000100011: out_v[345] = 10'b0010000101;
    16'b0010000101000010: out_v[345] = 10'b1100010011;
    16'b0110000001100011: out_v[345] = 10'b0010011111;
    16'b0110000001000010: out_v[345] = 10'b1101011011;
    16'b0010011101100011: out_v[345] = 10'b0010001101;
    16'b0010001001100011: out_v[345] = 10'b1010101011;
    16'b0010000001100011: out_v[345] = 10'b1001011011;
    16'b0110000001100010: out_v[345] = 10'b1010010011;
    16'b0010000101100011: out_v[345] = 10'b0110111110;
    16'b0010010100100011: out_v[345] = 10'b1111001011;
    16'b0010000101100010: out_v[345] = 10'b1001100110;
    16'b0000000100100010: out_v[345] = 10'b1101011101;
    16'b0000010101100010: out_v[345] = 10'b0010110110;
    16'b0010010101100011: out_v[345] = 10'b0011111101;
    16'b0010011101100000: out_v[345] = 10'b1011110111;
    16'b0000010101100011: out_v[345] = 10'b0010101111;
    16'b0010011101100001: out_v[345] = 10'b1000101111;
    16'b0010000001000010: out_v[345] = 10'b1010111111;
    16'b0110010001100011: out_v[345] = 10'b1011100111;
    16'b0010010101100010: out_v[345] = 10'b1011011111;
    16'b0000010100100011: out_v[345] = 10'b0000000011;
    16'b0000000001000010: out_v[345] = 10'b1001010101;
    16'b0010010100100010: out_v[345] = 10'b1011101111;
    16'b0010011101100010: out_v[345] = 10'b1011110110;
    16'b0110000101000010: out_v[345] = 10'b0010011011;
    16'b0000000100100011: out_v[345] = 10'b1001010001;
    16'b0000000001000000: out_v[345] = 10'b0111110000;
    16'b0000000101100010: out_v[345] = 10'b1011110110;
    16'b0110000101100011: out_v[345] = 10'b1001001011;
    16'b0110000001000001: out_v[345] = 10'b0001111001;
    16'b0010010001100011: out_v[345] = 10'b1011111100;
    16'b0000010000100011: out_v[345] = 10'b0110010111;
    16'b0010010000100011: out_v[345] = 10'b1110001100;
    16'b0000000001000011: out_v[345] = 10'b1001011010;
    16'b0000000000100011: out_v[345] = 10'b0110111001;
    16'b0110000011000000: out_v[345] = 10'b0100011100;
    16'b0010000011000000: out_v[345] = 10'b1100100111;
    16'b0000000010000010: out_v[345] = 10'b1011011001;
    16'b0110000010000000: out_v[345] = 10'b0000011101;
    16'b0000000010000000: out_v[345] = 10'b1001110010;
    16'b0000000010100010: out_v[345] = 10'b1011001011;
    16'b0000000011000000: out_v[345] = 10'b1101100011;
    16'b0010000010000000: out_v[345] = 10'b0101011011;
    16'b0100000011000000: out_v[345] = 10'b1011000011;
    16'b0010000010000010: out_v[345] = 10'b0101010010;
    16'b0000010010100010: out_v[345] = 10'b1011001011;
    16'b0000001010100010: out_v[345] = 10'b1110101111;
    16'b0010001010000000: out_v[345] = 10'b1001111111;
    16'b0110000011000001: out_v[345] = 10'b0011000111;
    16'b0000001010000000: out_v[345] = 10'b1000101111;
    16'b0000000011000001: out_v[345] = 10'b1001001010;
    16'b0000001010000010: out_v[345] = 10'b1001001101;
    16'b0010001011000000: out_v[345] = 10'b1110001100;
    16'b0010001010000010: out_v[345] = 10'b1010000110;
    16'b0110000010000010: out_v[345] = 10'b1011011001;
    16'b0110000011000010: out_v[345] = 10'b0010110001;
    16'b0010000010100010: out_v[345] = 10'b1110000011;
    16'b0010010010100011: out_v[345] = 10'b0000001110;
    16'b0010010011100010: out_v[345] = 10'b0011011001;
    16'b0000010010100000: out_v[345] = 10'b0110101001;
    16'b0110000011000011: out_v[345] = 10'b0011000111;
    16'b0000000010000011: out_v[345] = 10'b1110100101;
    16'b0010000010000011: out_v[345] = 10'b0010111010;
    16'b0000000000000010: out_v[345] = 10'b0101010110;
    16'b0110000011100001: out_v[345] = 10'b0100110110;
    16'b0000000010000001: out_v[345] = 10'b0111000110;
    16'b0110010011100001: out_v[345] = 10'b0001111011;
    16'b0110010001100001: out_v[345] = 10'b0011101011;
    16'b0110010011100011: out_v[345] = 10'b0100011111;
    16'b0110000011100000: out_v[345] = 10'b0101001100;
    16'b0010000011100001: out_v[345] = 10'b0011100011;
    16'b0010000000000001: out_v[345] = 10'b0110010100;
    16'b0010000000000011: out_v[345] = 10'b0010011101;
    16'b0010000011000001: out_v[345] = 10'b0111100000;
    16'b0010000011000010: out_v[345] = 10'b0010110001;
    16'b0010010010100001: out_v[345] = 10'b1100011111;
    16'b0000010000100010: out_v[345] = 10'b1001000101;
    16'b0000010010100001: out_v[345] = 10'b0100001101;
    16'b0010010010100010: out_v[345] = 10'b0010011010;
    16'b0110010001100010: out_v[345] = 10'b0101110110;
    16'b0000010000100001: out_v[345] = 10'b1100001111;
    16'b0000000010100001: out_v[345] = 10'b1101001010;
    16'b0000000000000001: out_v[345] = 10'b0000101111;
    16'b0010000010000001: out_v[345] = 10'b0000011101;
    16'b0110000011100011: out_v[345] = 10'b0101001110;
    16'b0010000011000011: out_v[345] = 10'b0111000111;
    16'b0010010011100001: out_v[345] = 10'b1111011111;
    16'b0000010010100011: out_v[345] = 10'b0011011101;
    16'b0010010001100001: out_v[345] = 10'b0101101111;
    16'b0000000000000011: out_v[345] = 10'b0000110101;
    16'b0110000001100001: out_v[345] = 10'b1001011001;
    16'b0110010011100000: out_v[345] = 10'b1111000100;
    16'b0010010011100011: out_v[345] = 10'b1100100111;
    16'b1000010010100001: out_v[345] = 10'b1000011101;
    16'b0110010011100010: out_v[345] = 10'b0011001001;
    16'b0000000010100011: out_v[345] = 10'b0011110100;
    16'b0010011010100010: out_v[345] = 10'b1101010101;
    16'b0110000011100010: out_v[345] = 10'b1110111011;
    16'b0000011010100000: out_v[345] = 10'b0011001111;
    16'b0000011010100010: out_v[345] = 10'b0100011110;
    16'b0010011011100000: out_v[345] = 10'b1010011001;
    16'b0010000011100010: out_v[345] = 10'b0111000001;
    16'b0010000000000010: out_v[345] = 10'b0101010011;
    16'b0010011011100010: out_v[345] = 10'b1011011011;
    16'b0000010110100010: out_v[345] = 10'b1100000100;
    16'b0000001010100000: out_v[345] = 10'b1101100101;
    16'b0000011011100010: out_v[345] = 10'b0010110001;
    16'b0010011010100000: out_v[345] = 10'b1011000101;
    16'b0000010011100010: out_v[345] = 10'b1101100001;
    16'b0010010001100010: out_v[345] = 10'b0001011110;
    16'b0010011011100011: out_v[345] = 10'b1000111010;
    16'b0000011000100010: out_v[345] = 10'b0001010001;
    16'b0000000000100010: out_v[345] = 10'b0001001111;
    16'b0000011110100010: out_v[345] = 10'b1101001010;
    16'b0010011111100010: out_v[345] = 10'b0011000011;
    16'b0000011010100011: out_v[345] = 10'b0110001000;
    16'b0010010000100010: out_v[345] = 10'b0001001110;
    16'b0010000111000001: out_v[345] = 10'b0111111011;
    16'b0000000100000001: out_v[345] = 10'b1000111000;
    16'b0000000111000001: out_v[345] = 10'b1100011001;
    16'b0000000110100000: out_v[345] = 10'b0001111011;
    16'b0000000101000001: out_v[345] = 10'b1001111110;
    16'b0000000110000010: out_v[345] = 10'b0110110000;
    16'b0000011111100010: out_v[345] = 10'b1001110101;
    16'b0000010110100011: out_v[345] = 10'b1111010000;
    16'b0000000110000000: out_v[345] = 10'b1010001111;
    16'b0010000110000010: out_v[345] = 10'b0011001100;
    16'b0000000010100000: out_v[345] = 10'b1001011001;
    16'b0000010100100001: out_v[345] = 10'b1001101010;
    16'b0010000110000001: out_v[345] = 10'b0110111100;
    16'b0000000110000011: out_v[345] = 10'b0101110010;
    16'b0000000110000001: out_v[345] = 10'b0110111011;
    16'b0000000111000010: out_v[345] = 10'b1111100111;
    16'b0000000111000000: out_v[345] = 10'b0011011101;
    16'b0000010111100011: out_v[345] = 10'b0010011011;
    16'b0000010110100001: out_v[345] = 10'b1110101010;
    16'b0000010110100000: out_v[345] = 10'b1001011111;
    16'b0000010111100010: out_v[345] = 10'b0100110011;
    16'b0000000001000001: out_v[345] = 10'b0100110011;
    16'b0000000100000011: out_v[345] = 10'b1001001011;
    16'b0000000100000000: out_v[345] = 10'b0110000101;
    16'b0000000101000011: out_v[345] = 10'b1100100110;
    16'b0000000011100000: out_v[345] = 10'b0010011001;
    16'b0010000100000001: out_v[345] = 10'b0111011011;
    16'b0000001111000010: out_v[345] = 10'b0101110110;
    16'b0000000111000011: out_v[345] = 10'b0110001010;
    16'b0010000110000000: out_v[345] = 10'b0111010011;
    16'b0010000111000010: out_v[345] = 10'b0010001110;
    16'b0000011111100011: out_v[345] = 10'b0001010101;
    16'b0000000011000011: out_v[345] = 10'b1010101110;
    16'b0000000000100001: out_v[345] = 10'b0010111001;
    16'b0000000000000000: out_v[345] = 10'b0010001001;
    16'b0010001011100010: out_v[345] = 10'b1110000001;
    16'b0010010111100010: out_v[345] = 10'b1011011010;
    16'b0010011111100000: out_v[345] = 10'b0110111111;
    16'b0000000011000010: out_v[345] = 10'b0100010011;
    16'b0010000111100010: out_v[345] = 10'b0101110001;
    16'b0000000011100010: out_v[345] = 10'b0111110111;
    16'b0000011111100000: out_v[345] = 10'b0111101110;
    16'b0010001111100010: out_v[345] = 10'b0011101001;
    16'b0110010111100010: out_v[345] = 10'b1010100101;
    16'b0000000110100010: out_v[345] = 10'b1100101010;
    16'b0110010010100010: out_v[345] = 10'b0100111001;
    16'b0000000111100010: out_v[345] = 10'b1111010100;
    16'b0110010110100010: out_v[345] = 10'b0110100110;
    16'b0110000010100011: out_v[345] = 10'b0111010110;
    16'b0010000010100011: out_v[345] = 10'b1101110000;
    16'b0110000000000011: out_v[345] = 10'b0011111000;
    16'b0110000000000010: out_v[345] = 10'b1111100010;
    16'b0110000111100011: out_v[345] = 10'b1011001010;
    16'b0110010110100011: out_v[345] = 10'b1001011010;
    16'b0110000010000011: out_v[345] = 10'b1100010101;
    16'b0110000110100011: out_v[345] = 10'b1111010010;
    16'b0110000000100011: out_v[345] = 10'b0101010010;
    16'b0110000000000001: out_v[345] = 10'b1011001010;
    16'b0110010111100011: out_v[345] = 10'b0111110011;
    16'b0010010110100011: out_v[345] = 10'b1111010011;
    16'b0000010110000011: out_v[345] = 10'b1111001111;
    16'b0110000010000001: out_v[345] = 10'b1011110101;
    16'b0110000010100010: out_v[345] = 10'b0110100100;
    16'b0000010000100000: out_v[345] = 10'b1011000010;
    16'b0000001100000010: out_v[345] = 10'b1000011100;
    16'b0000000100000010: out_v[345] = 10'b0111100000;
    16'b0000001000000010: out_v[345] = 10'b0011000011;
    16'b0000001000100010: out_v[345] = 10'b0110110100;
    16'b0000000000100000: out_v[345] = 10'b1110101010;
    16'b0000010011100000: out_v[345] = 10'b0111010001;
    16'b0000100100000000: out_v[345] = 10'b0010011110;
    16'b0000001100100010: out_v[345] = 10'b1101100000;
    16'b0000100000000000: out_v[345] = 10'b0111001101;
    16'b0000011100100010: out_v[345] = 10'b0111001101;
    16'b0000001110000010: out_v[345] = 10'b0000111011;
    16'b0000100000100000: out_v[345] = 10'b0101011111;
    16'b0000000100100000: out_v[345] = 10'b1010101000;
    16'b0000001110100010: out_v[345] = 10'b1111000001;
    16'b0000110000100000: out_v[345] = 10'b1101111101;
    16'b0000010100100000: out_v[345] = 10'b1011100010;
    16'b0000100100100000: out_v[345] = 10'b1111101011;
    16'b0000100110000000: out_v[345] = 10'b1101000111;
    16'b0000010001100000: out_v[345] = 10'b0011101000;
    16'b0010010110100010: out_v[345] = 10'b0110100101;
    16'b0010001011100011: out_v[345] = 10'b0110011110;
    16'b0010011110100010: out_v[345] = 10'b1011100100;
    16'b0010000011100011: out_v[345] = 10'b1100100010;
    16'b0010010111100011: out_v[345] = 10'b0110010010;
    16'b0000011110100000: out_v[345] = 10'b1011110010;
    16'b0010011011100001: out_v[345] = 10'b1010101110;
    16'b0010011111100001: out_v[345] = 10'b0101000000;
    16'b0010011111100011: out_v[345] = 10'b1110110110;
    16'b0000001111100010: out_v[345] = 10'b1111001101;
    16'b0000001011100010: out_v[345] = 10'b0101010111;
    16'b0000000111100000: out_v[345] = 10'b1011110011;
    16'b0000000110100011: out_v[345] = 10'b0010111010;
    16'b0000001110100011: out_v[345] = 10'b1100011110;
    16'b0000001111100011: out_v[345] = 10'b0011111101;
    16'b0000001011000011: out_v[345] = 10'b1011000111;
    16'b0000000111100011: out_v[345] = 10'b1110000111;
    16'b0000011110100011: out_v[345] = 10'b1101011101;
    16'b0000000100100001: out_v[345] = 10'b1100010011;
    16'b0000000110100001: out_v[345] = 10'b1000100111;
    default: out_v[345] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0101000010000000: out_v[346] = 10'b0100100000;
    16'b0101001010100101: out_v[346] = 10'b0100001011;
    16'b0101001010100001: out_v[346] = 10'b1011011110;
    16'b0100000010000100: out_v[346] = 10'b1111011001;
    16'b0100001010000101: out_v[346] = 10'b1110010110;
    16'b0100000010100101: out_v[346] = 10'b1111101010;
    16'b0100001000100001: out_v[346] = 10'b1010011101;
    16'b0000001010100001: out_v[346] = 10'b1000010111;
    16'b0001001010100001: out_v[346] = 10'b1001001011;
    16'b0101000010000100: out_v[346] = 10'b1111001001;
    16'b0100001010100001: out_v[346] = 10'b0000110111;
    16'b0101001010000001: out_v[346] = 10'b0111100001;
    16'b0100001010100101: out_v[346] = 10'b1110000001;
    16'b0100000010000000: out_v[346] = 10'b1000101011;
    16'b0101001010000101: out_v[346] = 10'b1100011111;
    16'b0101000010100001: out_v[346] = 10'b1001000010;
    16'b0100000010100001: out_v[346] = 10'b1111001001;
    16'b0100001000000101: out_v[346] = 10'b0101100101;
    16'b0101001010000100: out_v[346] = 10'b1110011010;
    16'b0100000010100000: out_v[346] = 10'b1111001100;
    16'b0100000000100001: out_v[346] = 10'b0000011101;
    16'b0111000010100001: out_v[346] = 10'b1011011111;
    16'b0101001010100000: out_v[346] = 10'b1010011111;
    16'b0100000010000101: out_v[346] = 10'b1010110101;
    16'b0001001010000000: out_v[346] = 10'b0000011111;
    16'b0000001010100101: out_v[346] = 10'b1001110010;
    16'b0000000010100101: out_v[346] = 10'b1011100101;
    16'b0101001000100001: out_v[346] = 10'b1011010001;
    16'b0101000010000101: out_v[346] = 10'b1001011011;
    16'b0101001000000100: out_v[346] = 10'b1010100010;
    16'b0100000010000001: out_v[346] = 10'b1000000110;
    16'b0001000010000000: out_v[346] = 10'b0100000010;
    16'b0101000010100101: out_v[346] = 10'b1110100010;
    16'b0101000000000100: out_v[346] = 10'b1000101011;
    16'b0100000000000100: out_v[346] = 10'b1110100000;
    16'b0101000010100000: out_v[346] = 10'b0110101011;
    16'b0101000010000001: out_v[346] = 10'b1100101010;
    16'b0101001010000000: out_v[346] = 10'b1010100101;
    16'b0100001010000001: out_v[346] = 10'b1010110010;
    16'b0111001010100001: out_v[346] = 10'b0111100110;
    16'b0000000010000100: out_v[346] = 10'b0011011110;
    16'b0101000000000000: out_v[346] = 10'b0101001010;
    16'b0100000000000000: out_v[346] = 10'b1001110010;
    16'b0000000000000100: out_v[346] = 10'b0011011101;
    16'b0000000000000000: out_v[346] = 10'b0111010100;
    16'b0001000000000100: out_v[346] = 10'b0110010100;
    16'b0000000010100100: out_v[346] = 10'b1001100011;
    16'b0001000000000000: out_v[346] = 10'b0010100011;
    16'b0110000000000100: out_v[346] = 10'b1100010100;
    16'b0110000010000100: out_v[346] = 10'b1100000111;
    16'b0000001010000100: out_v[346] = 10'b0110111010;
    16'b0100000000000101: out_v[346] = 10'b0100110100;
    16'b0010000010000100: out_v[346] = 10'b0001111100;
    16'b0110001000000100: out_v[346] = 10'b1001101110;
    16'b0110000000000000: out_v[346] = 10'b0010110100;
    16'b0000000010000101: out_v[346] = 10'b1000011000;
    16'b0110001000000101: out_v[346] = 10'b1110011010;
    16'b0001000010000100: out_v[346] = 10'b0101010011;
    16'b0110001010000101: out_v[346] = 10'b0010101111;
    16'b0111000010000100: out_v[346] = 10'b1001011111;
    16'b0000001000000000: out_v[346] = 10'b1011001101;
    16'b0110001010000100: out_v[346] = 10'b1101010010;
    16'b0111000000000100: out_v[346] = 10'b0011101110;
    16'b0010000000000100: out_v[346] = 10'b1000010010;
    16'b0110000010000101: out_v[346] = 10'b0000011100;
    16'b0100001010000100: out_v[346] = 10'b1100001100;
    16'b0000000010000001: out_v[346] = 10'b0000110111;
    16'b0100001000000100: out_v[346] = 10'b0100110111;
    16'b0110000000000101: out_v[346] = 10'b0110001111;
    16'b0000001000000100: out_v[346] = 10'b0011110100;
    16'b0000000010100001: out_v[346] = 10'b1101000001;
    16'b0110001000000000: out_v[346] = 10'b0010101011;
    16'b0100000000100000: out_v[346] = 10'b1100011110;
    16'b0000000010000000: out_v[346] = 10'b1100100101;
    16'b0100001000000000: out_v[346] = 10'b0011011010;
    16'b0000001010000000: out_v[346] = 10'b1110000011;
    16'b0100001010000000: out_v[346] = 10'b0110110001;
    16'b0000001010000101: out_v[346] = 10'b0011111011;
    16'b0101001000000000: out_v[346] = 10'b0010111101;
    16'b0001001010000100: out_v[346] = 10'b0100000011;
    16'b0111001000000100: out_v[346] = 10'b1010011111;
    16'b0001001000000000: out_v[346] = 10'b1010110110;
    16'b0101001010100100: out_v[346] = 10'b1001110001;
    16'b0100000010100100: out_v[346] = 10'b1011110000;
    16'b0111001010000100: out_v[346] = 10'b1100111000;
    16'b0001001000000100: out_v[346] = 10'b1100101001;
    16'b0101000010100100: out_v[346] = 10'b1001110110;
    16'b0001000000100000: out_v[346] = 10'b0110011011;
    16'b0000000000100000: out_v[346] = 10'b0010010110;
    16'b0001000010000001: out_v[346] = 10'b0101111110;
    16'b0001001010000101: out_v[346] = 10'b1010011011;
    16'b0000000000000101: out_v[346] = 10'b0010011101;
    16'b0000000000100001: out_v[346] = 10'b0100011011;
    16'b0001000010000101: out_v[346] = 10'b0100010111;
    16'b0101000000100001: out_v[346] = 10'b1111001111;
    16'b0001000010100001: out_v[346] = 10'b1111111111;
    16'b0000001010000001: out_v[346] = 10'b0000110011;
    16'b0001000000100001: out_v[346] = 10'b0010011001;
    16'b0000000000100100: out_v[346] = 10'b0010101000;
    16'b0000000010100000: out_v[346] = 10'b1101001000;
    16'b0111001000000000: out_v[346] = 10'b0011101110;
    16'b0000000000100101: out_v[346] = 10'b0011101000;
    16'b0001000010100100: out_v[346] = 10'b0000110001;
    16'b0101001000000001: out_v[346] = 10'b0101111010;
    16'b0101000000000001: out_v[346] = 10'b0010110010;
    16'b0100010000000000: out_v[346] = 10'b1010010010;
    16'b1100011000000000: out_v[346] = 10'b0001111111;
    16'b0000001000000001: out_v[346] = 10'b0111000111;
    16'b0100001000000001: out_v[346] = 10'b1011011010;
    16'b0000000000000001: out_v[346] = 10'b0011000000;
    16'b1100001000000001: out_v[346] = 10'b1111001010;
    16'b1100000000000000: out_v[346] = 10'b0011011001;
    16'b0000010000000000: out_v[346] = 10'b0010110010;
    16'b0100011000000000: out_v[346] = 10'b1111011010;
    16'b0000001000000101: out_v[346] = 10'b1010000011;
    16'b1100011000000001: out_v[346] = 10'b1111101110;
    16'b1000010000000000: out_v[346] = 10'b1111001010;
    16'b0100011000000001: out_v[346] = 10'b1111011010;
    16'b1100001000000000: out_v[346] = 10'b1010110111;
    16'b1100010000000000: out_v[346] = 10'b0110110101;
    16'b0001000010100101: out_v[346] = 10'b1011000100;
    16'b0001000000100100: out_v[346] = 10'b1110101111;
    16'b0100000000100100: out_v[346] = 10'b1111110111;
    16'b0101000000100100: out_v[346] = 10'b0000100111;
    16'b0101000000100000: out_v[346] = 10'b1100011111;
    default: out_v[346] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100111001110001: out_v[347] = 10'b1011011100;
    16'b0000111001010000: out_v[347] = 10'b0100101101;
    16'b0000110001110001: out_v[347] = 10'b1111010000;
    16'b0100111001010001: out_v[347] = 10'b1011011011;
    16'b0100101100100000: out_v[347] = 10'b1000111001;
    16'b0000110001010001: out_v[347] = 10'b1011100010;
    16'b0000100000000000: out_v[347] = 10'b0000111111;
    16'b0000111001010001: out_v[347] = 10'b1011010011;
    16'b0100111101110001: out_v[347] = 10'b1010011011;
    16'b0000100000000001: out_v[347] = 10'b1100011010;
    16'b0100111101110000: out_v[347] = 10'b1101000000;
    16'b0000001001010001: out_v[347] = 10'b1110011101;
    16'b0100011001010001: out_v[347] = 10'b0000101001;
    16'b0000100100000000: out_v[347] = 10'b0101000101;
    16'b0100111101010001: out_v[347] = 10'b0010101010;
    16'b0000111101110001: out_v[347] = 10'b1001001010;
    16'b0000101101010001: out_v[347] = 10'b1001010000;
    16'b0100111001100001: out_v[347] = 10'b0111000101;
    16'b0001110001010001: out_v[347] = 10'b1011010011;
    16'b0000110001010000: out_v[347] = 10'b0010110000;
    16'b0000111001110001: out_v[347] = 10'b0000101011;
    16'b0001110001010000: out_v[347] = 10'b0010001111;
    16'b0000010001010001: out_v[347] = 10'b0011001001;
    16'b0000101100000000: out_v[347] = 10'b0110101011;
    16'b0000011001010001: out_v[347] = 10'b0000011101;
    16'b0100101101110000: out_v[347] = 10'b1100010011;
    16'b0000111101010001: out_v[347] = 10'b0011101010;
    16'b0000101101110000: out_v[347] = 10'b0011100111;
    16'b0000111101010000: out_v[347] = 10'b1010110110;
    16'b0000010001010000: out_v[347] = 10'b1001011001;
    16'b0000000001010001: out_v[347] = 10'b0001111001;
    16'b0101111001010001: out_v[347] = 10'b1000010110;
    16'b0000111101110000: out_v[347] = 10'b0011111011;
    16'b0100101101110001: out_v[347] = 10'b1010110110;
    16'b0000101101010000: out_v[347] = 10'b0010101100;
    16'b0100111000100001: out_v[347] = 10'b0011010111;
    16'b0000110101010001: out_v[347] = 10'b0001001110;
    16'b0100101100000000: out_v[347] = 10'b1001010001;
    16'b0100111000000001: out_v[347] = 10'b0100000111;
    16'b0000011001010000: out_v[347] = 10'b1100010111;
    16'b0100100100000000: out_v[347] = 10'b0001101101;
    16'b0000110000000001: out_v[347] = 10'b1000100011;
    16'b0100100001110000: out_v[347] = 10'b0100110011;
    16'b0000010000000000: out_v[347] = 10'b1111000111;
    16'b0000110001000001: out_v[347] = 10'b0010111111;
    16'b0000010000000001: out_v[347] = 10'b1011000100;
    16'b0000000000000001: out_v[347] = 10'b0111100111;
    16'b0000100001010000: out_v[347] = 10'b1111100111;
    16'b0000100001010001: out_v[347] = 10'b0110001011;
    16'b0000010100000001: out_v[347] = 10'b0101010001;
    16'b0100000000000000: out_v[347] = 10'b0000111010;
    16'b0000000100000001: out_v[347] = 10'b0011011001;
    16'b0100000000010000: out_v[347] = 10'b0001111111;
    16'b0100001000100000: out_v[347] = 10'b1001111011;
    16'b0100100001010001: out_v[347] = 10'b1100110001;
    16'b0000000100000000: out_v[347] = 10'b1000010111;
    16'b0000110001000000: out_v[347] = 10'b1011101001;
    16'b0000100000010000: out_v[347] = 10'b0101010110;
    16'b0100100101110000: out_v[347] = 10'b1010110010;
    16'b0100100001010000: out_v[347] = 10'b0001101111;
    16'b0100100000100000: out_v[347] = 10'b1101011000;
    16'b0100000000100000: out_v[347] = 10'b1010010011;
    16'b0000100001000001: out_v[347] = 10'b0111010010;
    16'b0100100000110000: out_v[347] = 10'b0111011011;
    16'b0100100000010000: out_v[347] = 10'b1110011101;
    16'b0100100000000000: out_v[347] = 10'b1010111000;
    16'b0000010001000001: out_v[347] = 10'b0011110101;
    16'b0000100101010000: out_v[347] = 10'b1000011100;
    16'b0000100001000000: out_v[347] = 10'b1011001001;
    16'b0000110101000001: out_v[347] = 10'b1000110011;
    16'b0000010100000000: out_v[347] = 10'b1100010001;
    16'b0000110100000001: out_v[347] = 10'b1111101011;
    16'b0000000000000000: out_v[347] = 10'b1000001001;
    16'b0000010101000001: out_v[347] = 10'b0001111111;
    16'b0100110001110001: out_v[347] = 10'b0000011100;
    16'b0100001100100000: out_v[347] = 10'b1001110101;
    16'b0100100000000001: out_v[347] = 10'b0001111101;
    16'b0100001100100001: out_v[347] = 10'b1010111000;
    16'b0100101100100001: out_v[347] = 10'b0011100100;
    16'b0000001100100000: out_v[347] = 10'b0111011011;
    16'b0110101100100001: out_v[347] = 10'b0111011010;
    16'b0000101100100001: out_v[347] = 10'b1011100100;
    16'b0110100100100001: out_v[347] = 10'b1111011111;
    16'b0100110001010001: out_v[347] = 10'b1010100111;
    16'b0100101000100001: out_v[347] = 10'b1011000010;
    16'b0100101100110001: out_v[347] = 10'b1000011111;
    16'b0100100100100001: out_v[347] = 10'b0111100100;
    16'b0100001100000001: out_v[347] = 10'b1000011101;
    16'b0000001100100001: out_v[347] = 10'b0010011111;
    16'b0010101100100001: out_v[347] = 10'b1111000110;
    16'b0110101100000001: out_v[347] = 10'b0000010111;
    16'b0100100101110001: out_v[347] = 10'b0110101110;
    16'b0100100000100001: out_v[347] = 10'b1111011100;
    16'b0100000100100001: out_v[347] = 10'b0011110100;
    16'b0100001100000000: out_v[347] = 10'b0000011110;
    16'b0000101100000001: out_v[347] = 10'b1110010111;
    16'b0000100100100001: out_v[347] = 10'b1001100011;
    16'b0100110101110001: out_v[347] = 10'b0010110111;
    16'b0100001000000001: out_v[347] = 10'b1000101011;
    16'b0100101000000001: out_v[347] = 10'b1010010101;
    16'b0110100100000001: out_v[347] = 10'b1010110100;
    16'b0000101101110001: out_v[347] = 10'b0101010000;
    16'b0110001100100001: out_v[347] = 10'b0011110110;
    16'b0110111100100001: out_v[347] = 10'b1011001110;
    16'b0100101100000001: out_v[347] = 10'b1111001100;
    16'b0000110101110001: out_v[347] = 10'b1001100111;
    16'b0100000100000001: out_v[347] = 10'b1100010010;
    16'b0100100100110001: out_v[347] = 10'b1101000010;
    16'b0100100100000001: out_v[347] = 10'b1000110111;
    16'b0100000100000000: out_v[347] = 10'b1010101101;
    16'b0100001000100001: out_v[347] = 10'b1001111100;
    16'b0100000100100000: out_v[347] = 10'b1011101110;
    16'b0000000001110001: out_v[347] = 10'b1011101010;
    16'b0000100101110001: out_v[347] = 10'b0101111000;
    16'b0000010101110000: out_v[347] = 10'b0101000111;
    16'b0000010101010001: out_v[347] = 10'b0011100110;
    16'b0000110101110000: out_v[347] = 10'b1010100011;
    16'b0000110000100001: out_v[347] = 10'b0100101010;
    16'b0000010101010000: out_v[347] = 10'b0001111100;
    16'b0000100101010001: out_v[347] = 10'b0111001111;
    16'b0000100100100000: out_v[347] = 10'b1011011000;
    16'b0000010001110001: out_v[347] = 10'b0000111010;
    16'b0000011001110001: out_v[347] = 10'b0111101010;
    16'b0010110000100001: out_v[347] = 10'b0111011011;
    16'b0000010101110001: out_v[347] = 10'b1001101010;
    16'b0010110000000001: out_v[347] = 10'b0010011001;
    16'b0000011101110001: out_v[347] = 10'b1011000111;
    16'b0000000101010001: out_v[347] = 10'b1011111000;
    16'b0000110001110000: out_v[347] = 10'b0100011110;
    16'b0000001100000000: out_v[347] = 10'b0100100111;
    16'b0000101001110000: out_v[347] = 10'b0001010101;
    16'b0000000100100000: out_v[347] = 10'b1001101101;
    16'b0001001100100000: out_v[347] = 10'b1001111111;
    16'b0100011101100000: out_v[347] = 10'b1100010110;
    16'b0000100101110000: out_v[347] = 10'b1010000001;
    16'b0000011100100000: out_v[347] = 10'b1011001010;
    16'b0000010101100000: out_v[347] = 10'b0011010010;
    16'b0000001000100000: out_v[347] = 10'b1110010010;
    16'b0000101100110000: out_v[347] = 10'b1000000111;
    16'b0100011100100000: out_v[347] = 10'b1000010100;
    16'b0000010100100000: out_v[347] = 10'b0111010010;
    16'b0000001100000001: out_v[347] = 10'b1000111010;
    16'b0101001100100000: out_v[347] = 10'b0011111011;
    16'b0001001000100000: out_v[347] = 10'b1010010100;
    16'b0000101100100000: out_v[347] = 10'b0001010111;
    16'b0000100001110000: out_v[347] = 10'b1101011101;
    16'b0001000100100000: out_v[347] = 10'b0011100111;
    16'b0000011100000000: out_v[347] = 10'b0010100010;
    16'b0000111101100000: out_v[347] = 10'b0010110101;
    16'b0000011101100000: out_v[347] = 10'b0111101110;
    16'b0100011100000000: out_v[347] = 10'b0011110010;
    16'b0100111101100000: out_v[347] = 10'b0101010110;
    16'b0000110101010000: out_v[347] = 10'b0000111111;
    16'b0000011101010000: out_v[347] = 10'b0101111111;
    16'b0000000001010000: out_v[347] = 10'b1001100011;
    16'b0000100100010000: out_v[347] = 10'b1111010010;
    16'b0000000101010000: out_v[347] = 10'b0011101110;
    16'b0000110100000000: out_v[347] = 10'b0110100001;
    16'b0000010001110000: out_v[347] = 10'b1101110101;
    16'b0100111100000001: out_v[347] = 10'b1011001000;
    16'b0110101100100000: out_v[347] = 10'b1110000011;
    16'b0100111100100001: out_v[347] = 10'b0111100101;
    16'b0100111100000000: out_v[347] = 10'b0001000110;
    16'b0100110100000001: out_v[347] = 10'b1000001010;
    16'b0110001000100000: out_v[347] = 10'b1100000100;
    16'b0100101000100000: out_v[347] = 10'b0111101011;
    16'b0100111000100000: out_v[347] = 10'b0111010101;
    16'b0110001100100000: out_v[347] = 10'b1111101011;
    16'b0100110100000000: out_v[347] = 10'b1011010111;
    16'b0100110000000001: out_v[347] = 10'b0000111111;
    16'b0110101000100000: out_v[347] = 10'b0000111011;
    16'b0100111000000000: out_v[347] = 10'b1100100011;
    16'b0100101000000000: out_v[347] = 10'b0011111000;
    16'b0110101000100001: out_v[347] = 10'b1011111111;
    16'b0110111000100000: out_v[347] = 10'b1011110110;
    16'b0001100101110000: out_v[347] = 10'b0011001011;
    16'b0001000000000000: out_v[347] = 10'b0110110000;
    16'b0001110101110000: out_v[347] = 10'b1010001011;
    16'b0000110101100000: out_v[347] = 10'b0001110110;
    16'b0001000000101000: out_v[347] = 10'b0011111001;
    16'b0001010100100000: out_v[347] = 10'b0111111011;
    16'b0000100100110000: out_v[347] = 10'b1001100001;
    16'b0001010101100000: out_v[347] = 10'b1000001111;
    16'b0000100000110000: out_v[347] = 10'b1110010000;
    16'b0000010101000000: out_v[347] = 10'b1010001001;
    16'b0001110101100000: out_v[347] = 10'b1101010010;
    16'b0000000000100000: out_v[347] = 10'b1010100101;
    16'b0001000000100000: out_v[347] = 10'b0011010101;
    16'b0001010101110000: out_v[347] = 10'b0110101011;
    16'b0100100100110000: out_v[347] = 10'b0011010010;
    16'b0100001101110001: out_v[347] = 10'b0111010011;
    16'b0100010101110001: out_v[347] = 10'b0111110010;
    16'b0100000101110001: out_v[347] = 10'b0111000010;
    16'b0100110101110000: out_v[347] = 10'b0100000111;
    16'b0100010001110001: out_v[347] = 10'b1001011110;
    16'b0100100001110001: out_v[347] = 10'b0101000001;
    16'b0100111001110000: out_v[347] = 10'b0010101011;
    16'b0100110101010001: out_v[347] = 10'b1000100001;
    16'b0100010101010001: out_v[347] = 10'b0111000001;
    16'b0100010101110000: out_v[347] = 10'b1111010001;
    16'b0100101001110001: out_v[347] = 10'b0001011000;
    16'b0100110001110000: out_v[347] = 10'b0111011101;
    16'b0100011101110000: out_v[347] = 10'b0001101011;
    16'b0100011001110001: out_v[347] = 10'b0110100010;
    16'b0100000001110001: out_v[347] = 10'b0011010101;
    16'b0100001001110001: out_v[347] = 10'b0101010111;
    16'b0100100101010001: out_v[347] = 10'b1101100110;
    16'b0100011101110001: out_v[347] = 10'b0101110001;
    16'b0100101001110000: out_v[347] = 10'b1110100100;
    16'b0100010001110000: out_v[347] = 10'b0111000101;
    16'b0000110101100001: out_v[347] = 10'b0110010101;
    16'b0100011101010001: out_v[347] = 10'b0100100110;
    16'b0000011101110000: out_v[347] = 10'b0011011100;
    16'b0101001000100000: out_v[347] = 10'b1100001111;
    default: out_v[347] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000100100001: out_v[348] = 10'b1100001011;
    16'b0000100101110000: out_v[348] = 10'b1011010111;
    16'b0000100011110000: out_v[348] = 10'b1111111110;
    16'b0000100101110001: out_v[348] = 10'b1000011001;
    16'b0000000101100000: out_v[348] = 10'b1011011011;
    16'b0000000101110001: out_v[348] = 10'b0000100110;
    16'b0000000011110000: out_v[348] = 10'b0100011011;
    16'b0000100001110001: out_v[348] = 10'b0111101110;
    16'b0000000001110000: out_v[348] = 10'b1000100110;
    16'b0000100100110000: out_v[348] = 10'b1011011011;
    16'b0000100101100001: out_v[348] = 10'b1100011110;
    16'b0000100100110001: out_v[348] = 10'b0100000101;
    16'b0000100101010000: out_v[348] = 10'b1001110110;
    16'b1001100101110001: out_v[348] = 10'b0101101010;
    16'b0000100100010000: out_v[348] = 10'b0011000110;
    16'b0000100110110000: out_v[348] = 10'b0100101111;
    16'b0000000100110000: out_v[348] = 10'b0011001011;
    16'b0000100001010000: out_v[348] = 10'b0011010001;
    16'b0000100100100001: out_v[348] = 10'b0001001010;
    16'b0000100111110001: out_v[348] = 10'b0011111100;
    16'b0000000001100001: out_v[348] = 10'b0100001111;
    16'b0000100101100000: out_v[348] = 10'b1000110100;
    16'b0000100001110000: out_v[348] = 10'b1111011010;
    16'b0000100111110000: out_v[348] = 10'b0011000011;
    16'b0000100101010001: out_v[348] = 10'b0111001001;
    16'b0000000101100001: out_v[348] = 10'b0100011011;
    16'b0000000111110000: out_v[348] = 10'b0111001111;
    16'b0000000101110000: out_v[348] = 10'b1001001011;
    16'b0000100001010001: out_v[348] = 10'b1101011011;
    16'b0000000001010000: out_v[348] = 10'b1011001011;
    16'b0000000111110001: out_v[348] = 10'b0111111110;
    16'b0000100100100000: out_v[348] = 10'b1011110111;
    16'b0000100000110000: out_v[348] = 10'b1010111111;
    16'b0001100101110001: out_v[348] = 10'b1010001111;
    16'b1001100001000000: out_v[348] = 10'b1000101010;
    16'b1001000001000000: out_v[348] = 10'b0111000111;
    16'b1001000000100000: out_v[348] = 10'b1000001001;
    16'b0000000001100000: out_v[348] = 10'b1010111011;
    16'b0000000000100000: out_v[348] = 10'b0010101010;
    16'b0000000100000000: out_v[348] = 10'b0011111011;
    16'b0001000001000000: out_v[348] = 10'b0010110100;
    16'b0000000101000000: out_v[348] = 10'b0011101100;
    16'b1001100000000000: out_v[348] = 10'b1000011011;
    16'b1001100101000000: out_v[348] = 10'b0110011011;
    16'b0001000000100000: out_v[348] = 10'b0001001111;
    16'b1001000101000000: out_v[348] = 10'b1110100101;
    16'b1001000001100000: out_v[348] = 10'b1111010000;
    16'b0001000101000000: out_v[348] = 10'b0011100101;
    16'b0001000100100000: out_v[348] = 10'b0110110101;
    16'b1001000101100000: out_v[348] = 10'b1110110110;
    16'b0001000101100000: out_v[348] = 10'b0101011101;
    16'b0000000100100000: out_v[348] = 10'b0010110011;
    16'b0000000001000000: out_v[348] = 10'b0111100010;
    16'b1001000100100000: out_v[348] = 10'b1010001111;
    16'b0000000000000000: out_v[348] = 10'b1000000111;
    16'b0001000001100000: out_v[348] = 10'b1100000010;
    16'b1001000100000000: out_v[348] = 10'b0100010111;
    16'b0001000100000000: out_v[348] = 10'b0111100111;
    16'b1001100101100000: out_v[348] = 10'b1001011111;
    16'b1001100101010000: out_v[348] = 10'b0111101000;
    16'b1001100101110000: out_v[348] = 10'b0001000100;
    16'b0000000101000001: out_v[348] = 10'b0101000110;
    16'b1001000011100000: out_v[348] = 10'b1100010100;
    16'b1001100101010001: out_v[348] = 10'b0111011110;
    16'b1001100100000000: out_v[348] = 10'b1010001000;
    16'b0001100101000000: out_v[348] = 10'b0110100101;
    16'b0000000001110001: out_v[348] = 10'b1100110110;
    16'b1001000101110000: out_v[348] = 10'b0011011100;
    16'b1001100101100001: out_v[348] = 10'b0000100010;
    16'b0000000101010001: out_v[348] = 10'b1110100110;
    16'b0000000100110001: out_v[348] = 10'b1110110010;
    16'b1001000100110000: out_v[348] = 10'b0000111111;
    16'b1001000001110000: out_v[348] = 10'b0111011010;
    16'b1001000000110000: out_v[348] = 10'b0110100111;
    16'b1001100111100000: out_v[348] = 10'b0111100110;
    16'b1001000100010000: out_v[348] = 10'b0100110101;
    16'b0000100101000001: out_v[348] = 10'b0110010101;
    16'b1001000111100000: out_v[348] = 10'b0100001110;
    16'b0000100100010001: out_v[348] = 10'b1010100111;
    16'b1001000101010000: out_v[348] = 10'b0100110111;
    16'b0001100101100001: out_v[348] = 10'b0001110111;
    16'b1001000101110001: out_v[348] = 10'b1101001110;
    16'b1001100110100001: out_v[348] = 10'b0010110010;
    16'b0001100100000000: out_v[348] = 10'b0110111000;
    16'b0000100100000000: out_v[348] = 10'b1010111110;
    16'b1001100101000001: out_v[348] = 10'b1100011000;
    16'b1001100000100000: out_v[348] = 10'b0110000100;
    16'b1001100100100000: out_v[348] = 10'b1011010011;
    16'b1001100100000001: out_v[348] = 10'b1111001001;
    16'b1001100100100001: out_v[348] = 10'b1011100110;
    16'b1001100001100001: out_v[348] = 10'b0001110110;
    16'b0001100100100000: out_v[348] = 10'b0110001110;
    16'b1001100110100000: out_v[348] = 10'b0101010010;
    16'b1001000000100001: out_v[348] = 10'b1011101010;
    16'b1001000001100001: out_v[348] = 10'b0011010101;
    16'b1001100000100001: out_v[348] = 10'b0010010001;
    16'b1001000010100000: out_v[348] = 10'b1011011001;
    16'b1001100100110000: out_v[348] = 10'b1101010011;
    16'b1001100100110001: out_v[348] = 10'b0111100000;
    16'b1001000101100001: out_v[348] = 10'b1011101010;
    16'b0001100101100000: out_v[348] = 10'b0101011100;
    16'b1001100001100000: out_v[348] = 10'b0111011001;
    16'b1001000100000001: out_v[348] = 10'b0011110101;
    16'b1001000001010000: out_v[348] = 10'b0000111000;
    16'b1001000000000000: out_v[348] = 10'b0001111001;
    16'b0000000000100001: out_v[348] = 10'b1011000111;
    16'b1001000001000001: out_v[348] = 10'b1001101000;
    16'b1001000010000000: out_v[348] = 10'b0011001101;
    16'b1001000001110001: out_v[348] = 10'b0000101111;
    16'b1001000010010001: out_v[348] = 10'b1010100111;
    16'b0001000001100001: out_v[348] = 10'b0100100011;
    16'b0000000000000001: out_v[348] = 10'b1101011100;
    16'b0000000001000001: out_v[348] = 10'b1111001100;
    16'b1001000010000001: out_v[348] = 10'b0011010100;
    16'b0001000001010001: out_v[348] = 10'b1111110110;
    16'b0000000000010001: out_v[348] = 10'b1010110000;
    16'b1001000000010001: out_v[348] = 10'b0001010110;
    16'b0000000010000001: out_v[348] = 10'b0011011001;
    16'b0001000000000001: out_v[348] = 10'b1101101011;
    16'b1001000000000001: out_v[348] = 10'b0110111011;
    16'b0001000001000001: out_v[348] = 10'b0011001111;
    16'b0000000000110001: out_v[348] = 10'b1011010010;
    16'b0001000000000000: out_v[348] = 10'b1001110110;
    16'b0001000010000001: out_v[348] = 10'b1001101111;
    16'b0000000010010001: out_v[348] = 10'b0110111010;
    16'b0000000001010001: out_v[348] = 10'b0011110011;
    16'b1001000000010000: out_v[348] = 10'b1111100111;
    16'b0001000000100001: out_v[348] = 10'b1001011110;
    16'b1001000110000001: out_v[348] = 10'b1001110111;
    16'b1001000001010001: out_v[348] = 10'b1011111001;
    16'b1001000110010001: out_v[348] = 10'b0111011011;
    16'b0001000000010001: out_v[348] = 10'b0000011100;
    16'b1001000000110001: out_v[348] = 10'b1010110010;
    16'b0000100001000000: out_v[348] = 10'b1000111001;
    16'b0000100000100000: out_v[348] = 10'b1101100101;
    16'b0000100000000000: out_v[348] = 10'b1011100110;
    16'b0000100001100000: out_v[348] = 10'b0010100100;
    16'b1001000100100001: out_v[348] = 10'b1110100111;
    16'b0000101001000000: out_v[348] = 10'b0111111001;
    16'b1001000111100001: out_v[348] = 10'b1011100000;
    16'b0001100001000000: out_v[348] = 10'b1011110001;
    16'b0000101000100000: out_v[348] = 10'b1111010110;
    16'b0000101100100000: out_v[348] = 10'b1000001110;
    16'b0001000101100001: out_v[348] = 10'b1111100111;
    16'b1001000011010001: out_v[348] = 10'b1010111011;
    16'b0001000101110001: out_v[348] = 10'b0110100111;
    16'b1001000011010000: out_v[348] = 10'b1011001010;
    16'b0000000101010000: out_v[348] = 10'b1101000100;
    16'b1001000101000001: out_v[348] = 10'b1001111100;
    16'b1001000101010001: out_v[348] = 10'b1110101010;
    16'b0000000011010001: out_v[348] = 10'b0011110010;
    16'b0000000011000001: out_v[348] = 10'b1101001110;
    16'b1001000011000000: out_v[348] = 10'b1100100110;
    16'b0000000010100001: out_v[348] = 10'b1010010000;
    16'b1001000010100001: out_v[348] = 10'b1000000111;
    16'b0000000011100001: out_v[348] = 10'b0100001011;
    16'b1001000011000001: out_v[348] = 10'b0111101011;
    16'b0000100001000001: out_v[348] = 10'b1101011100;
    16'b0001100001100001: out_v[348] = 10'b1011100000;
    16'b0000000010000000: out_v[348] = 10'b0111110110;
    16'b1001000011100001: out_v[348] = 10'b0100101111;
    16'b0000100001100001: out_v[348] = 10'b0111001110;
    16'b0001000010100001: out_v[348] = 10'b1000001111;
    16'b1001100001000001: out_v[348] = 10'b1010101010;
    16'b0001000011100001: out_v[348] = 10'b1101010101;
    16'b0001000011000001: out_v[348] = 10'b0101101001;
    16'b0000100011100001: out_v[348] = 10'b0100010110;
    16'b0001100100100001: out_v[348] = 10'b1000010110;
    16'b0000000010110001: out_v[348] = 10'b0111100010;
    16'b1001000010110001: out_v[348] = 10'b1000101010;
    16'b0001000000110001: out_v[348] = 10'b0101000010;
    16'b1011000000100000: out_v[348] = 10'b1011000111;
    default: out_v[348] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001000100000001: out_v[349] = 10'b0111011001;
    16'b0101011100000001: out_v[349] = 10'b1001010101;
    16'b0101001100000001: out_v[349] = 10'b1000101001;
    16'b1101011100000001: out_v[349] = 10'b0100110100;
    16'b0001001100000001: out_v[349] = 10'b0100111101;
    16'b0101001000000001: out_v[349] = 10'b0001011100;
    16'b1100001000000000: out_v[349] = 10'b1001000000;
    16'b1100001100000001: out_v[349] = 10'b1010110101;
    16'b1000000100000001: out_v[349] = 10'b1100001001;
    16'b1101001000000001: out_v[349] = 10'b0001010101;
    16'b0000000100000001: out_v[349] = 10'b1111000111;
    16'b0101001000000000: out_v[349] = 10'b1011100100;
    16'b0001001000000001: out_v[349] = 10'b0001111000;
    16'b1101001100000001: out_v[349] = 10'b0000110111;
    16'b0101001100000000: out_v[349] = 10'b0010011000;
    16'b1100001000000001: out_v[349] = 10'b1010110100;
    16'b0001000000000001: out_v[349] = 10'b1001101100;
    16'b1000001100000001: out_v[349] = 10'b1110111011;
    16'b0100001100000001: out_v[349] = 10'b1001101101;
    16'b1000010100000001: out_v[349] = 10'b0111010011;
    16'b0100011100000001: out_v[349] = 10'b0100001011;
    16'b1001000100000001: out_v[349] = 10'b1111100010;
    16'b0101011100000000: out_v[349] = 10'b1000110011;
    16'b1000011100000001: out_v[349] = 10'b1110001010;
    16'b1000000000000001: out_v[349] = 10'b1000001110;
    16'b0001001000000000: out_v[349] = 10'b0100110101;
    16'b1100101000000001: out_v[349] = 10'b0011000001;
    16'b0001011100000001: out_v[349] = 10'b1001010110;
    16'b1100011100000001: out_v[349] = 10'b0000001111;
    16'b0000001100000001: out_v[349] = 10'b1110000101;
    16'b0001000000000000: out_v[349] = 10'b0000010101;
    16'b0101011000000001: out_v[349] = 10'b0110001010;
    16'b1000001000000001: out_v[349] = 10'b0000100111;
    16'b0100001000000001: out_v[349] = 10'b0010010110;
    16'b1000000100000000: out_v[349] = 10'b0110100111;
    16'b0000001000000000: out_v[349] = 10'b1001101101;
    16'b0000000000000000: out_v[349] = 10'b0110111101;
    16'b0100001000000000: out_v[349] = 10'b0001010110;
    16'b0000000000000001: out_v[349] = 10'b0110100011;
    16'b0000010000000000: out_v[349] = 10'b1011010010;
    16'b0000001000000001: out_v[349] = 10'b1100101001;
    16'b0000000100000000: out_v[349] = 10'b0000010010;
    16'b0000010000000001: out_v[349] = 10'b1011011001;
    16'b1000000000000000: out_v[349] = 10'b0001100101;
    16'b1001000000000000: out_v[349] = 10'b1000001011;
    16'b1001000000000001: out_v[349] = 10'b0000101100;
    16'b0001010000000001: out_v[349] = 10'b0111110110;
    16'b0100011000000001: out_v[349] = 10'b0001011100;
    16'b0000011100000001: out_v[349] = 10'b0010111111;
    16'b1000001000000000: out_v[349] = 10'b1101101111;
    16'b1001001000000001: out_v[349] = 10'b1010110000;
    16'b1100011000000001: out_v[349] = 10'b0110010001;
    16'b1001001000000000: out_v[349] = 10'b1101001011;
    16'b1101001000000000: out_v[349] = 10'b0111001110;
    16'b0000010100000001: out_v[349] = 10'b1100001100;
    16'b0000011000000001: out_v[349] = 10'b0000111111;
    16'b0001010100000001: out_v[349] = 10'b0111101000;
    16'b0001000100000000: out_v[349] = 10'b1001010010;
    16'b1001000100000000: out_v[349] = 10'b0111010000;
    16'b1001011100000001: out_v[349] = 10'b0101010110;
    16'b1001010100000001: out_v[349] = 10'b0111101010;
    16'b1001001100000001: out_v[349] = 10'b1010110110;
    16'b0100001100000000: out_v[349] = 10'b0100110011;
    16'b0001001100000000: out_v[349] = 10'b0101110110;
    16'b0000001100000000: out_v[349] = 10'b0111010000;
    16'b0110001000000000: out_v[349] = 10'b1001110001;
    16'b0010001000000000: out_v[349] = 10'b1001001111;
    16'b0111001000000000: out_v[349] = 10'b0111010000;
    16'b0110001000000001: out_v[349] = 10'b1111000001;
    16'b0101101000000000: out_v[349] = 10'b1010101001;
    16'b0001100000000000: out_v[349] = 10'b1010001101;
    16'b0100011100000000: out_v[349] = 10'b0101100110;
    16'b0000010100000000: out_v[349] = 10'b1100000100;
    16'b0011000000000010: out_v[349] = 10'b0111110011;
    16'b0011000000000000: out_v[349] = 10'b1001101111;
    16'b0010000000000000: out_v[349] = 10'b1000101100;
    16'b0111001000000010: out_v[349] = 10'b1101011011;
    16'b0100001100001000: out_v[349] = 10'b0011100111;
    16'b0011001000000000: out_v[349] = 10'b0010011110;
    16'b0111001000000001: out_v[349] = 10'b1101000111;
    16'b0010000100000001: out_v[349] = 10'b0101010111;
    16'b0110001100000001: out_v[349] = 10'b0101011111;
    16'b0010001000000001: out_v[349] = 10'b1110100011;
    16'b0011000000000001: out_v[349] = 10'b1001101010;
    16'b0010000000000001: out_v[349] = 10'b0001101100;
    16'b0001100000000001: out_v[349] = 10'b1000001001;
    16'b0011001000000001: out_v[349] = 10'b1111001000;
    default: out_v[349] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0110100000000110: out_v[350] = 10'b0110000111;
    16'b1010000000100110: out_v[350] = 10'b0101101110;
    16'b1010000000100100: out_v[350] = 10'b0010010001;
    16'b1010000000110100: out_v[350] = 10'b1011010101;
    16'b1000100000100010: out_v[350] = 10'b0100111001;
    16'b1000000000100000: out_v[350] = 10'b0000001011;
    16'b1000000000100010: out_v[350] = 10'b0100100011;
    16'b1000100000100000: out_v[350] = 10'b0100110101;
    16'b0010000000010100: out_v[350] = 10'b0001101010;
    16'b1110100000000110: out_v[350] = 10'b1111010001;
    16'b1111100000100110: out_v[350] = 10'b1000010011;
    16'b0010000000000110: out_v[350] = 10'b1010101100;
    16'b0010100000000100: out_v[350] = 10'b0010011001;
    16'b0010000001010100: out_v[350] = 10'b0000100011;
    16'b1010000000000110: out_v[350] = 10'b1011110110;
    16'b1110100000100110: out_v[350] = 10'b1010011001;
    16'b1000000000110000: out_v[350] = 10'b0001011011;
    16'b0010100000110100: out_v[350] = 10'b0101011001;
    16'b0010000000110100: out_v[350] = 10'b0110110101;
    16'b0010000001000100: out_v[350] = 10'b0100100111;
    16'b0010000000100100: out_v[350] = 10'b1001110110;
    16'b1100100000100010: out_v[350] = 10'b0101000001;
    16'b0000000000100000: out_v[350] = 10'b0101000011;
    16'b1000100000110000: out_v[350] = 10'b0011110010;
    16'b1010100000100110: out_v[350] = 10'b1011111110;
    16'b0010000000000100: out_v[350] = 10'b0110011011;
    16'b0010100001110100: out_v[350] = 10'b0010001111;
    16'b0110100000010110: out_v[350] = 10'b1110000011;
    16'b0010100000010100: out_v[350] = 10'b1001011101;
    16'b1010100000100100: out_v[350] = 10'b0111001000;
    16'b0010100001010100: out_v[350] = 10'b1111011111;
    16'b1010100000110100: out_v[350] = 10'b0111011010;
    16'b1100000000100010: out_v[350] = 10'b1111101011;
    16'b1010100000110110: out_v[350] = 10'b0011111110;
    16'b1110100000110110: out_v[350] = 10'b0100000011;
    16'b0010000001110100: out_v[350] = 10'b1011110100;
    16'b0010100000000110: out_v[350] = 10'b0011111110;
    16'b1101100000100010: out_v[350] = 10'b0101100001;
    16'b1010000000110110: out_v[350] = 10'b1101000110;
    16'b0110100000110110: out_v[350] = 10'b0001100111;
    16'b0100100000100000: out_v[350] = 10'b0000101111;
    16'b0000000000000000: out_v[350] = 10'b0111000111;
    16'b0100100000000000: out_v[350] = 10'b0000010110;
    16'b1000000000000000: out_v[350] = 10'b0001001111;
    16'b0000100000000000: out_v[350] = 10'b1011111010;
    16'b1010000000000100: out_v[350] = 10'b0111101101;
    16'b1000000000010000: out_v[350] = 10'b1001000011;
    16'b0100000000100000: out_v[350] = 10'b1010100010;
    16'b0101100000100000: out_v[350] = 10'b0011100010;
    16'b1111000000100100: out_v[350] = 10'b1010100010;
    16'b0100100000000010: out_v[350] = 10'b0011010010;
    16'b1101100000100000: out_v[350] = 10'b0100000100;
    16'b1011000000100100: out_v[350] = 10'b0111010011;
    16'b1011000000110100: out_v[350] = 10'b0111111010;
    16'b0100100000100010: out_v[350] = 10'b0111000000;
    16'b0110000000100100: out_v[350] = 10'b0011101001;
    16'b0101100000000000: out_v[350] = 10'b1010001110;
    16'b0100000000000000: out_v[350] = 10'b1110110111;
    16'b1010000000010100: out_v[350] = 10'b0101111001;
    16'b1001000000010000: out_v[350] = 10'b0001000111;
    16'b0000100000100000: out_v[350] = 10'b1100111011;
    16'b1100100000100000: out_v[350] = 10'b0100010101;
    16'b1110000000100100: out_v[350] = 10'b0100011001;
    16'b0110100001110100: out_v[350] = 10'b0011110011;
    16'b1101100001110000: out_v[350] = 10'b0011001011;
    16'b1101000000110010: out_v[350] = 10'b1011101011;
    16'b1001100000110000: out_v[350] = 10'b0111100000;
    16'b0111100001110100: out_v[350] = 10'b0111010011;
    16'b1100100001110000: out_v[350] = 10'b0110011101;
    16'b1100100000110000: out_v[350] = 10'b0101001110;
    16'b1101100000110000: out_v[350] = 10'b0100001010;
    16'b0110100001010100: out_v[350] = 10'b1111010111;
    16'b1001100000100000: out_v[350] = 10'b0101111100;
    16'b1101100000110010: out_v[350] = 10'b1001011100;
    16'b1001100001110000: out_v[350] = 10'b1111000101;
    16'b1101000000110000: out_v[350] = 10'b0010111001;
    16'b1101100000000000: out_v[350] = 10'b0110001011;
    16'b1100100000110010: out_v[350] = 10'b1110000110;
    16'b1100000000110000: out_v[350] = 10'b1100000110;
    16'b1100100000000000: out_v[350] = 10'b0101100101;
    16'b1001000001110000: out_v[350] = 10'b0000010101;
    16'b1101000000100000: out_v[350] = 10'b1101100100;
    16'b0101100000010000: out_v[350] = 10'b0111100011;
    16'b1111100000110100: out_v[350] = 10'b1100010110;
    16'b1101100001010000: out_v[350] = 10'b0110011010;
    16'b1101000001110000: out_v[350] = 10'b0111110011;
    16'b0110100000010100: out_v[350] = 10'b0011010101;
    16'b0101100000000010: out_v[350] = 10'b0010010100;
    16'b1111100001110100: out_v[350] = 10'b1011110100;
    16'b1101100001110010: out_v[350] = 10'b1010001111;
    16'b1101100000010000: out_v[350] = 10'b0100111011;
    16'b1001000000110010: out_v[350] = 10'b0010110111;
    16'b1001000000110000: out_v[350] = 10'b1111110010;
    16'b1100100000010000: out_v[350] = 10'b1101100100;
    16'b1100100001110010: out_v[350] = 10'b0101010110;
    16'b0101100000110000: out_v[350] = 10'b1011010101;
    16'b1101100001100000: out_v[350] = 10'b0010111011;
    16'b1100000000100000: out_v[350] = 10'b0101100100;
    16'b0100100000110000: out_v[350] = 10'b1011011101;
    16'b0010000000010110: out_v[350] = 10'b1001000100;
    16'b0011000000010110: out_v[350] = 10'b1111000101;
    16'b0011000001010110: out_v[350] = 10'b1111101110;
    16'b0010000000110110: out_v[350] = 10'b0111100101;
    16'b0111000000000100: out_v[350] = 10'b1001001000;
    16'b0110000000000110: out_v[350] = 10'b0010101101;
    16'b0011000001010100: out_v[350] = 10'b0011011001;
    16'b1001000000100010: out_v[350] = 10'b0011100110;
    16'b1111000000100110: out_v[350] = 10'b1000011110;
    16'b1011000000110110: out_v[350] = 10'b0101010111;
    16'b0011000000000100: out_v[350] = 10'b1101011000;
    16'b0110000001010110: out_v[350] = 10'b0011111000;
    16'b0011000000000110: out_v[350] = 10'b0001100110;
    16'b1000000000110010: out_v[350] = 10'b1010010110;
    16'b1101000000100010: out_v[350] = 10'b0000111000;
    16'b0110000000010110: out_v[350] = 10'b1000101010;
    16'b0010000001110110: out_v[350] = 10'b1011000000;
    16'b0010000001010110: out_v[350] = 10'b0110000110;
    16'b1111000000010110: out_v[350] = 10'b0010011100;
    16'b0111000000010110: out_v[350] = 10'b1011101111;
    16'b1000001000100010: out_v[350] = 10'b1111001010;
    16'b0111000001010110: out_v[350] = 10'b0011111111;
    16'b1011000000000110: out_v[350] = 10'b1100010010;
    16'b1111000000110110: out_v[350] = 10'b0010111011;
    16'b1011000000010110: out_v[350] = 10'b1101001001;
    16'b1111000000000110: out_v[350] = 10'b1000000101;
    16'b0011000000110110: out_v[350] = 10'b1111000111;
    16'b0111000000010100: out_v[350] = 10'b0111111001;
    16'b0011000000010100: out_v[350] = 10'b0111111001;
    16'b1110000000000110: out_v[350] = 10'b0010101110;
    16'b1010000000010110: out_v[350] = 10'b0101011100;
    16'b0111000000000110: out_v[350] = 10'b1000101111;
    16'b1011000000010100: out_v[350] = 10'b0101100111;
    16'b1001000000100000: out_v[350] = 10'b1001011100;
    16'b1101100000000010: out_v[350] = 10'b0011111111;
    16'b0101100000100010: out_v[350] = 10'b1101001010;
    16'b1011000000100110: out_v[350] = 10'b1111000101;
    16'b1101000000000000: out_v[350] = 10'b1100101001;
    16'b0101000000000010: out_v[350] = 10'b0000110100;
    16'b1001000000000010: out_v[350] = 10'b0101011100;
    16'b0101000000100010: out_v[350] = 10'b1001010001;
    16'b1111000000000100: out_v[350] = 10'b1111010001;
    16'b0001000000000010: out_v[350] = 10'b0110110101;
    16'b0101000000000000: out_v[350] = 10'b1100010001;
    16'b1101000000000010: out_v[350] = 10'b0010100111;
    16'b0101000001000000: out_v[350] = 10'b0001111111;
    16'b0101100001000000: out_v[350] = 10'b0000011000;
    16'b0101000001000010: out_v[350] = 10'b0011111011;
    16'b0101000000010000: out_v[350] = 10'b0100101000;
    16'b1111100000000110: out_v[350] = 10'b0011010000;
    16'b0001000000100010: out_v[350] = 10'b1011010001;
    16'b1111000000010100: out_v[350] = 10'b1010100010;
    16'b1111100000000100: out_v[350] = 10'b0110001011;
    16'b1111100000100100: out_v[350] = 10'b0010011010;
    16'b0101000000100000: out_v[350] = 10'b1011110001;
    16'b1001100000100010: out_v[350] = 10'b1110101011;
    16'b1110000000100110: out_v[350] = 10'b0110100111;
    16'b0110000000000100: out_v[350] = 10'b1001101010;
    16'b0010000001000110: out_v[350] = 10'b1100110100;
    16'b1110000000000100: out_v[350] = 10'b1001101100;
    16'b0100000000100010: out_v[350] = 10'b0100110110;
    16'b0011000001000110: out_v[350] = 10'b0011100111;
    16'b1001100000110010: out_v[350] = 10'b0010011110;
    16'b0100100000110010: out_v[350] = 10'b1111010011;
    16'b1001000010100000: out_v[350] = 10'b0101111110;
    16'b0001000010100000: out_v[350] = 10'b0001110111;
    16'b1011000000000100: out_v[350] = 10'b0100101111;
    16'b0000000001001000: out_v[350] = 10'b0110010110;
    16'b1001000010100010: out_v[350] = 10'b0111001011;
    16'b0000000000001000: out_v[350] = 10'b0111000100;
    16'b0001000000100000: out_v[350] = 10'b1111001010;
    16'b1001000000000000: out_v[350] = 10'b1111100011;
    16'b1000000010100000: out_v[350] = 10'b0110111001;
    16'b1011000010100100: out_v[350] = 10'b0110000110;
    16'b1001000000001000: out_v[350] = 10'b0111101001;
    16'b1010000010100100: out_v[350] = 10'b0111110110;
    16'b0001100000100000: out_v[350] = 10'b0111010011;
    16'b1110100000010110: out_v[350] = 10'b1110001011;
    16'b0111100000000110: out_v[350] = 10'b0111000110;
    16'b0110100000100110: out_v[350] = 10'b0100011000;
    16'b0111100000100110: out_v[350] = 10'b0111010000;
    16'b0111100000010110: out_v[350] = 10'b0101000010;
    16'b0111100000110110: out_v[350] = 10'b0110110110;
    16'b1110100000100100: out_v[350] = 10'b1111100001;
    16'b1111100000110110: out_v[350] = 10'b1011111001;
    16'b0111100001110110: out_v[350] = 10'b1110001010;
    16'b0111100001010110: out_v[350] = 10'b0110000000;
    16'b1111100000010100: out_v[350] = 10'b0110100111;
    16'b0111100000010100: out_v[350] = 10'b0111110110;
    16'b1111100000010110: out_v[350] = 10'b0110001111;
    16'b0111100000000100: out_v[350] = 10'b0111101100;
    16'b0110100001010110: out_v[350] = 10'b1110000111;
    16'b1110100000000100: out_v[350] = 10'b1100010100;
    16'b0011000000100110: out_v[350] = 10'b0110110101;
    16'b1011100000000110: out_v[350] = 10'b1000011011;
    16'b0111100001000110: out_v[350] = 10'b0111000110;
    16'b1101000010100000: out_v[350] = 10'b1000110001;
    16'b1101000010100010: out_v[350] = 10'b1111001111;
    16'b0101000000001000: out_v[350] = 10'b1001101011;
    16'b0100000000001000: out_v[350] = 10'b1100100101;
    16'b0001100000000000: out_v[350] = 10'b1001001011;
    16'b1101000000001000: out_v[350] = 10'b1110100111;
    16'b0101100000001000: out_v[350] = 10'b1001100011;
    16'b0100000001000000: out_v[350] = 10'b1000001011;
    default: out_v[350] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1001010000000000: out_v[351] = 10'b0001111001;
    16'b1011100000000010: out_v[351] = 10'b0111101111;
    16'b1011100000100010: out_v[351] = 10'b0011111110;
    16'b1011100001100010: out_v[351] = 10'b1000010111;
    16'b1011010000000010: out_v[351] = 10'b0010011111;
    16'b1010100001100010: out_v[351] = 10'b1100111011;
    16'b0011000000000000: out_v[351] = 10'b0111001110;
    16'b1001100001000010: out_v[351] = 10'b1000100111;
    16'b0010100001100010: out_v[351] = 10'b1111011110;
    16'b1011010000000000: out_v[351] = 10'b0110111001;
    16'b1011100001000010: out_v[351] = 10'b0101101100;
    16'b0011100000000010: out_v[351] = 10'b0110001011;
    16'b1001000000000000: out_v[351] = 10'b1100110010;
    16'b1001000000000010: out_v[351] = 10'b0101011001;
    16'b1011000000000010: out_v[351] = 10'b0101000001;
    16'b1011000000000000: out_v[351] = 10'b1111001011;
    16'b1001010000000010: out_v[351] = 10'b0010111111;
    16'b0011000000000010: out_v[351] = 10'b0001001001;
    16'b1011100000000000: out_v[351] = 10'b0100100001;
    16'b1000100000100000: out_v[351] = 10'b1110011011;
    16'b1001100000100010: out_v[351] = 10'b0111100011;
    16'b1010100001100000: out_v[351] = 10'b1011000111;
    16'b1011000000100010: out_v[351] = 10'b0011000101;
    16'b0001100000000010: out_v[351] = 10'b0110101111;
    16'b1001100000000000: out_v[351] = 10'b0000011101;
    16'b1000100001100000: out_v[351] = 10'b0100011001;
    16'b0011100001000010: out_v[351] = 10'b0101100010;
    16'b1001100000000010: out_v[351] = 10'b1010111111;
    16'b1000100001100010: out_v[351] = 10'b1110000001;
    16'b1010100001000010: out_v[351] = 10'b1111100011;
    16'b1011110001100010: out_v[351] = 10'b1010111011;
    16'b0011010000000010: out_v[351] = 10'b0001011010;
    16'b1000010000000000: out_v[351] = 10'b0110000110;
    16'b0000010000000000: out_v[351] = 10'b0101010101;
    16'b0001000000000000: out_v[351] = 10'b0110100111;
    16'b0010100001000010: out_v[351] = 10'b0111110010;
    16'b1011110000000010: out_v[351] = 10'b1110010011;
    16'b0001000000000010: out_v[351] = 10'b0101000111;
    16'b0100000000000000: out_v[351] = 10'b0101000001;
    16'b0000000000000000: out_v[351] = 10'b0000111011;
    16'b1000110000000000: out_v[351] = 10'b1111101001;
    16'b1001110000000000: out_v[351] = 10'b1011000110;
    16'b1000000000000000: out_v[351] = 10'b1000101100;
    16'b1001110000010000: out_v[351] = 10'b0000111111;
    16'b1000100000000000: out_v[351] = 10'b0010011010;
    16'b0001010000000000: out_v[351] = 10'b0010110101;
    16'b1000110000010000: out_v[351] = 10'b0010010101;
    16'b1001110001000010: out_v[351] = 10'b0111110110;
    16'b1001110000000010: out_v[351] = 10'b0101011100;
    16'b0001110001010000: out_v[351] = 10'b1110010101;
    16'b1001110001010000: out_v[351] = 10'b0011100110;
    16'b1001110001000000: out_v[351] = 10'b0011011100;
    16'b0001100000000000: out_v[351] = 10'b1101110101;
    16'b0001110000000000: out_v[351] = 10'b0110000110;
    16'b1001100001000000: out_v[351] = 10'b0111001111;
    16'b1000110001000000: out_v[351] = 10'b1010100011;
    16'b0001010000000010: out_v[351] = 10'b1100001110;
    16'b0000110000000000: out_v[351] = 10'b1011101011;
    16'b0001110001000010: out_v[351] = 10'b0111001110;
    16'b0001110001000000: out_v[351] = 10'b1101001101;
    16'b0001010000010000: out_v[351] = 10'b1010100111;
    16'b0001110000010000: out_v[351] = 10'b1010011101;
    16'b1001010000010000: out_v[351] = 10'b1000101101;
    16'b1001100000010000: out_v[351] = 10'b0011000100;
    16'b0000010000010000: out_v[351] = 10'b0011000001;
    16'b1000100001000010: out_v[351] = 10'b0111011100;
    16'b1000100001000000: out_v[351] = 10'b0010001010;
    16'b0000100001000000: out_v[351] = 10'b0000111000;
    16'b1010100001000000: out_v[351] = 10'b1011111001;
    16'b0000000000000010: out_v[351] = 10'b0010101010;
    16'b0010000000000000: out_v[351] = 10'b0000110110;
    16'b1100000000000000: out_v[351] = 10'b0011110111;
    16'b0000100000000010: out_v[351] = 10'b1011110110;
    16'b0000000000000110: out_v[351] = 10'b1010011011;
    16'b0010100000000000: out_v[351] = 10'b0011110100;
    16'b0000100000000000: out_v[351] = 10'b0000111010;
    16'b1010100000000000: out_v[351] = 10'b1111001000;
    16'b1000000000000010: out_v[351] = 10'b0011001100;
    16'b1000100000000010: out_v[351] = 10'b1011011000;
    16'b1010000000000000: out_v[351] = 10'b1011001110;
    16'b1000000010000000: out_v[351] = 10'b1101000000;
    16'b0010000000000010: out_v[351] = 10'b0010110110;
    16'b0000000000000100: out_v[351] = 10'b0001001101;
    16'b1000100001010000: out_v[351] = 10'b1011001111;
    16'b0000100001000010: out_v[351] = 10'b1011001110;
    16'b0011010000000000: out_v[351] = 10'b1001100000;
    16'b1001010000100000: out_v[351] = 10'b1001100111;
    16'b0110000000000000: out_v[351] = 10'b0011011101;
    16'b1010000000000010: out_v[351] = 10'b1001100110;
    16'b1011010000100000: out_v[351] = 10'b0001011011;
    16'b0010010000000010: out_v[351] = 10'b1111001011;
    16'b1010010000000000: out_v[351] = 10'b0100110000;
    16'b0010000000100010: out_v[351] = 10'b0010011110;
    16'b0010000000100000: out_v[351] = 10'b0010111110;
    16'b0010010000000000: out_v[351] = 10'b1100110010;
    16'b1010000000100010: out_v[351] = 10'b1001110110;
    16'b1011010000100010: out_v[351] = 10'b1110111011;
    16'b1010000000100000: out_v[351] = 10'b0001111110;
    16'b0011010000100010: out_v[351] = 10'b1100011011;
    16'b1110000000000000: out_v[351] = 10'b0000110111;
    16'b0011010000100000: out_v[351] = 10'b0111101011;
    16'b1010010000000010: out_v[351] = 10'b1101010110;
    16'b1110010000000000: out_v[351] = 10'b1000110111;
    16'b0010100001000000: out_v[351] = 10'b1100100110;
    16'b0010100000000010: out_v[351] = 10'b1001110100;
    16'b0011010000010000: out_v[351] = 10'b0011011010;
    16'b0011010000010010: out_v[351] = 10'b0001001101;
    16'b0001010000010010: out_v[351] = 10'b1010100100;
    16'b0000010000000010: out_v[351] = 10'b1011100111;
    16'b0011000000010000: out_v[351] = 10'b1101010000;
    16'b0001000000010010: out_v[351] = 10'b1011000110;
    16'b0011110000010010: out_v[351] = 10'b1101110110;
    16'b0011000000010010: out_v[351] = 10'b1111000010;
    16'b0011100000010010: out_v[351] = 10'b0111111000;
    16'b0001000000010000: out_v[351] = 10'b0111100000;
    16'b0000010000010010: out_v[351] = 10'b1011010000;
    16'b0000000000010000: out_v[351] = 10'b1000100010;
    16'b1110000000100000: out_v[351] = 10'b0011101111;
    16'b1000000010000010: out_v[351] = 10'b1110010011;
    16'b1100000000000100: out_v[351] = 10'b1001001110;
    16'b0100000000000100: out_v[351] = 10'b1001111011;
    16'b1000010010000000: out_v[351] = 10'b1010111011;
    16'b1010000010000000: out_v[351] = 10'b0111100010;
    16'b1000000000000100: out_v[351] = 10'b1000101010;
    16'b1101010000000000: out_v[351] = 10'b0011111001;
    16'b1100000000000110: out_v[351] = 10'b0111110000;
    16'b1100010000000000: out_v[351] = 10'b0101010111;
    16'b0100000000000110: out_v[351] = 10'b0110010111;
    16'b0100010000000000: out_v[351] = 10'b1101001001;
    16'b0110010000000000: out_v[351] = 10'b1101101000;
    16'b1111010000000000: out_v[351] = 10'b1000100101;
    16'b1001010000100010: out_v[351] = 10'b1100010001;
    16'b0111010000000000: out_v[351] = 10'b1101100011;
    16'b0001010000100000: out_v[351] = 10'b1101010011;
    default: out_v[351] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001000010100000: out_v[352] = 10'b0100100101;
    16'b0001000011100001: out_v[352] = 10'b0011110110;
    16'b0001000010101000: out_v[352] = 10'b0111001001;
    16'b0001000010100001: out_v[352] = 10'b1010010010;
    16'b0000000010000001: out_v[352] = 10'b1000000001;
    16'b0000000000000000: out_v[352] = 10'b0001110010;
    16'b0000000010000011: out_v[352] = 10'b0111100110;
    16'b0000000010001000: out_v[352] = 10'b1010111110;
    16'b0001000011100000: out_v[352] = 10'b1101011011;
    16'b0001000011101000: out_v[352] = 10'b0101011010;
    16'b0001000001100000: out_v[352] = 10'b1110010010;
    16'b0001000000100000: out_v[352] = 10'b1100010111;
    16'b0000000010000000: out_v[352] = 10'b0001001010;
    16'b0001001010100000: out_v[352] = 10'b1100011110;
    16'b0001000010100010: out_v[352] = 10'b0011010100;
    16'b0001001010100010: out_v[352] = 10'b0100000111;
    16'b0000001010000001: out_v[352] = 10'b0101000001;
    16'b0000000001000001: out_v[352] = 10'b0001110011;
    16'b0001000010101010: out_v[352] = 10'b0100011100;
    16'b0000000011000000: out_v[352] = 10'b0110111011;
    16'b0001001000100000: out_v[352] = 10'b1100010001;
    16'b0000000011000001: out_v[352] = 10'b0110100111;
    16'b0001001010100001: out_v[352] = 10'b1011000111;
    16'b0001000010101001: out_v[352] = 10'b1011011000;
    16'b0001000011100010: out_v[352] = 10'b1101110101;
    16'b0000000000001000: out_v[352] = 10'b0110010111;
    16'b0001000000100010: out_v[352] = 10'b1111000101;
    16'b0000000011001000: out_v[352] = 10'b1101000110;
    16'b0000010000000000: out_v[352] = 10'b0010011001;
    16'b0000000001000000: out_v[352] = 10'b0010011110;
    16'b0000000000000010: out_v[352] = 10'b0100100100;
    16'b0000000001001000: out_v[352] = 10'b0001011000;
    16'b0000000010001010: out_v[352] = 10'b0000001110;
    16'b0000000000001010: out_v[352] = 10'b0010110100;
    16'b0000000010000010: out_v[352] = 10'b0000101110;
    16'b0000001000001000: out_v[352] = 10'b0100011110;
    16'b0001000000101000: out_v[352] = 10'b0011110100;
    16'b0000000001000010: out_v[352] = 10'b1001011111;
    16'b0000000011001010: out_v[352] = 10'b1100100100;
    16'b0000000011000010: out_v[352] = 10'b1011001010;
    16'b0000010000001000: out_v[352] = 10'b1111101111;
    16'b0000010001000000: out_v[352] = 10'b0000111011;
    16'b0001000011101010: out_v[352] = 10'b1011111011;
    16'b0000000001001010: out_v[352] = 10'b0110111011;
    16'b0001000001101010: out_v[352] = 10'b1111001010;
    16'b0001000001101000: out_v[352] = 10'b1000001011;
    16'b0001001000101000: out_v[352] = 10'b1111100100;
    16'b0001000000101010: out_v[352] = 10'b0000010011;
    16'b0001000011101001: out_v[352] = 10'b0011011100;
    16'b0001000000100001: out_v[352] = 10'b0000111100;
    16'b0001010000101000: out_v[352] = 10'b1010101101;
    16'b0001000001101001: out_v[352] = 10'b0101011011;
    16'b0001000000101001: out_v[352] = 10'b1110001011;
    16'b0000000000000001: out_v[352] = 10'b0000101101;
    16'b0000010011000000: out_v[352] = 10'b0101010011;
    16'b0000000010001001: out_v[352] = 10'b1011110111;
    16'b0001010000100000: out_v[352] = 10'b1110001010;
    16'b0001011000100000: out_v[352] = 10'b1011110110;
    16'b0001010001101000: out_v[352] = 10'b1011001001;
    16'b0100001000001000: out_v[352] = 10'b1111010011;
    16'b0001001001101000: out_v[352] = 10'b1011110100;
    16'b0000011000001000: out_v[352] = 10'b0011110011;
    16'b0001000001100001: out_v[352] = 10'b0011111010;
    16'b0001011000101000: out_v[352] = 10'b1100001011;
    16'b0001001001100000: out_v[352] = 10'b1011110001;
    16'b0001011001101000: out_v[352] = 10'b0110111011;
    16'b0001011000101100: out_v[352] = 10'b0001011111;
    16'b0101001000101000: out_v[352] = 10'b1111001110;
    16'b0001010011101000: out_v[352] = 10'b0001110111;
    16'b0001010011101001: out_v[352] = 10'b0101110111;
    16'b0100000000001000: out_v[352] = 10'b1110000001;
    default: out_v[352] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000010000001100: out_v[353] = 10'b1001111101;
    16'b0000010000010100: out_v[353] = 10'b1100110010;
    16'b0100010100011100: out_v[353] = 10'b1111000111;
    16'b0000010000011100: out_v[353] = 10'b1101011100;
    16'b0000010000001000: out_v[353] = 10'b1011000100;
    16'b0000000000010100: out_v[353] = 10'b0000110101;
    16'b0011110000001100: out_v[353] = 10'b0111001000;
    16'b0100010100001100: out_v[353] = 10'b0010100101;
    16'b0000010100001100: out_v[353] = 10'b1010100011;
    16'b0000000000000100: out_v[353] = 10'b0010010011;
    16'b0000000000001100: out_v[353] = 10'b0011010110;
    16'b0000110000001100: out_v[353] = 10'b1010010001;
    16'b0000010100011100: out_v[353] = 10'b1101001001;
    16'b0000000000011100: out_v[353] = 10'b0110010010;
    16'b0100000100000100: out_v[353] = 10'b1110011101;
    16'b0100010110001100: out_v[353] = 10'b0000001011;
    16'b0000010000011000: out_v[353] = 10'b1111111001;
    16'b0000110000000100: out_v[353] = 10'b1110110111;
    16'b0000010000000100: out_v[353] = 10'b1000111001;
    16'b0000000100000100: out_v[353] = 10'b1110100100;
    16'b0000100000001100: out_v[353] = 10'b0111011101;
    16'b0000010000101100: out_v[353] = 10'b1000001011;
    16'b0000110000011100: out_v[353] = 10'b1101111101;
    16'b0011110000011100: out_v[353] = 10'b0011110011;
    16'b0011110000001000: out_v[353] = 10'b0000101110;
    16'b0011100000001100: out_v[353] = 10'b0100110000;
    16'b0011000000000100: out_v[353] = 10'b0101111101;
    16'b0011100000000000: out_v[353] = 10'b0000111101;
    16'b0011000000000000: out_v[353] = 10'b1001000110;
    16'b0011100000000100: out_v[353] = 10'b1000011101;
    16'b0011000000001000: out_v[353] = 10'b1100001011;
    16'b0010000000000100: out_v[353] = 10'b0000100011;
    16'b0010000000000000: out_v[353] = 10'b1000100111;
    16'b0011100000001000: out_v[353] = 10'b1000010101;
    16'b0011010000001000: out_v[353] = 10'b1101000111;
    16'b0000000000001000: out_v[353] = 10'b0011000111;
    16'b0000000000000000: out_v[353] = 10'b1000010010;
    16'b0011000000001100: out_v[353] = 10'b0110001101;
    16'b0011110000101100: out_v[353] = 10'b1011000000;
    16'b0011110100001100: out_v[353] = 10'b1001100100;
    16'b0000010000101000: out_v[353] = 10'b1011101110;
    16'b0011110100101100: out_v[353] = 10'b0011111010;
    16'b0000000100001100: out_v[353] = 10'b0011110110;
    16'b0011110000000000: out_v[353] = 10'b0100100111;
    16'b0111110100001000: out_v[353] = 10'b1000000110;
    16'b0111110100001100: out_v[353] = 10'b0100001000;
    16'b0000000000101000: out_v[353] = 10'b1100111010;
    16'b0000110000101000: out_v[353] = 10'b1110010111;
    16'b0000010100101000: out_v[353] = 10'b1100011100;
    16'b0011110000101000: out_v[353] = 10'b1000110101;
    16'b0011110100001000: out_v[353] = 10'b1011101100;
    16'b0100000100001100: out_v[353] = 10'b1000110101;
    16'b0011010000001100: out_v[353] = 10'b1100100101;
    16'b0011110100101000: out_v[353] = 10'b0011000111;
    16'b0000010100001000: out_v[353] = 10'b1110110010;
    16'b0011100000101000: out_v[353] = 10'b0110001100;
    16'b0111110110001100: out_v[353] = 10'b1101101111;
    16'b0000110000001000: out_v[353] = 10'b0110110001;
    16'b0100010100001000: out_v[353] = 10'b1000000111;
    16'b0010110000001000: out_v[353] = 10'b1101011010;
    16'b0011110000011000: out_v[353] = 10'b1010110011;
    16'b0000010100101100: out_v[353] = 10'b1110100101;
    16'b0000010000000000: out_v[353] = 10'b1100010110;
    16'b0111100100000100: out_v[353] = 10'b0001101010;
    16'b0011100110000100: out_v[353] = 10'b1011011000;
    16'b0011100100000100: out_v[353] = 10'b0010100101;
    16'b0011100100000000: out_v[353] = 10'b1010011010;
    16'b0111100110000100: out_v[353] = 10'b0110101011;
    16'b0011110000000100: out_v[353] = 10'b0111010000;
    16'b0011100110001100: out_v[353] = 10'b0000101001;
    16'b0011110110001100: out_v[353] = 10'b1010001111;
    16'b0111100110000000: out_v[353] = 10'b0011001111;
    16'b0011100100001100: out_v[353] = 10'b1101001001;
    16'b0111100100000000: out_v[353] = 10'b1000000011;
    16'b0111100110001100: out_v[353] = 10'b0100111000;
    16'b0011110100000100: out_v[353] = 10'b0100001000;
    16'b0111100100001100: out_v[353] = 10'b1111001010;
    16'b0011100110000000: out_v[353] = 10'b0001011010;
    16'b0000100100000100: out_v[353] = 10'b0010001100;
    16'b0000100000000100: out_v[353] = 10'b0110111110;
    16'b0010100000000100: out_v[353] = 10'b1010101010;
    16'b0100000100000000: out_v[353] = 10'b1011101001;
    16'b0011100000010100: out_v[353] = 10'b1001100010;
    16'b0011100000011100: out_v[353] = 10'b1100011011;
    16'b0111100010000000: out_v[353] = 10'b0001010111;
    16'b0111100000000000: out_v[353] = 10'b1100011001;
    16'b0010100000000000: out_v[353] = 10'b1000111101;
    16'b0000100100000000: out_v[353] = 10'b0011010000;
    16'b0000000100000000: out_v[353] = 10'b0011001101;
    16'b0011100000011000: out_v[353] = 10'b1100000100;
    16'b0000100000000000: out_v[353] = 10'b0100110001;
    16'b0000000000010000: out_v[353] = 10'b0000111111;
    16'b0000100000011100: out_v[353] = 10'b1011110000;
    16'b0000110000011000: out_v[353] = 10'b0111101111;
    16'b0000100000010100: out_v[353] = 10'b0011001011;
    16'b0011010000101000: out_v[353] = 10'b0101011011;
    16'b0010110000001100: out_v[353] = 10'b1011001001;
    16'b0000100000100000: out_v[353] = 10'b1011000110;
    16'b0011100000100000: out_v[353] = 10'b1111000101;
    16'b0000100000001000: out_v[353] = 10'b0101000001;
    16'b0000000000100000: out_v[353] = 10'b0001001110;
    16'b0011100000101100: out_v[353] = 10'b1011100110;
    16'b0100000000000000: out_v[353] = 10'b0111000000;
    16'b0100000110000000: out_v[353] = 10'b0111000010;
    16'b0100000110000100: out_v[353] = 10'b1100100110;
    16'b0100000000000100: out_v[353] = 10'b0001110100;
    16'b0100000010000100: out_v[353] = 10'b1101100010;
    16'b0100000000000010: out_v[353] = 10'b0011110010;
    16'b0000000000011000: out_v[353] = 10'b0011010101;
    16'b0100000000010100: out_v[353] = 10'b0001101101;
    16'b0100000010000000: out_v[353] = 10'b0111110011;
    16'b0000000110000100: out_v[353] = 10'b1110010011;
    16'b0000000100001000: out_v[353] = 10'b1010100010;
    16'b0011110000010100: out_v[353] = 10'b0111010010;
    16'b0111110100011100: out_v[353] = 10'b0001000010;
    16'b0011110100011100: out_v[353] = 10'b1000011011;
    default: out_v[353] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000001000010: out_v[354] = 10'b0010010000;
    16'b0000000000100010: out_v[354] = 10'b1101001001;
    16'b0100000001100000: out_v[354] = 10'b0110100101;
    16'b0100000001100010: out_v[354] = 10'b0010101101;
    16'b0000000000000010: out_v[354] = 10'b1011100011;
    16'b0100000001000000: out_v[354] = 10'b0000101101;
    16'b0100000000000000: out_v[354] = 10'b0011010010;
    16'b0000000001001010: out_v[354] = 10'b1110100011;
    16'b0000000000100000: out_v[354] = 10'b0010110010;
    16'b0100000000100010: out_v[354] = 10'b0010000001;
    16'b0100000001001010: out_v[354] = 10'b1010111011;
    16'b0100000001000010: out_v[354] = 10'b1010111010;
    16'b0000000001100000: out_v[354] = 10'b1010110000;
    16'b0000000000000000: out_v[354] = 10'b0001110010;
    16'b0100000001101010: out_v[354] = 10'b0101011000;
    16'b0000000001100010: out_v[354] = 10'b0010011000;
    16'b0000000001001000: out_v[354] = 10'b1001110010;
    16'b0000000001000000: out_v[354] = 10'b1110011000;
    16'b0100000000000010: out_v[354] = 10'b0011010001;
    16'b0100000001001000: out_v[354] = 10'b1001010101;
    16'b0100000000100000: out_v[354] = 10'b1001011101;
    16'b0000000000001000: out_v[354] = 10'b1000001100;
    16'b0000000010001000: out_v[354] = 10'b0011100100;
    16'b0100000011001010: out_v[354] = 10'b1010100111;
    16'b0000000001101000: out_v[354] = 10'b1101010001;
    16'b0000000001101010: out_v[354] = 10'b0111011000;
    16'b0100000000001010: out_v[354] = 10'b0100001011;
    16'b0000000010001010: out_v[354] = 10'b0101011011;
    16'b0000000000001010: out_v[354] = 10'b0010011010;
    16'b0000000011001010: out_v[354] = 10'b1000010111;
    16'b0100000000001000: out_v[354] = 10'b1100011100;
    16'b0000000011000000: out_v[354] = 10'b1001100101;
    16'b0000000011000010: out_v[354] = 10'b1111100110;
    16'b0000000000101010: out_v[354] = 10'b1101000110;
    16'b0000000011001000: out_v[354] = 10'b0011000111;
    16'b0000000011101010: out_v[354] = 10'b0110110011;
    16'b0000000000101000: out_v[354] = 10'b1101010101;
    16'b0100000000101000: out_v[354] = 10'b0000101111;
    16'b0100000000101010: out_v[354] = 10'b0111100111;
    16'b0100000011000000: out_v[354] = 10'b1010101101;
    16'b0100000011000010: out_v[354] = 10'b0100100011;
    default: out_v[354] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100100000000000: out_v[355] = 10'b0001110110;
    16'b0000100010000000: out_v[355] = 10'b1010010101;
    16'b0100100010000000: out_v[355] = 10'b1100011011;
    16'b0000100000000000: out_v[355] = 10'b0001110001;
    16'b0101000010000000: out_v[355] = 10'b0101011010;
    16'b0000000010000100: out_v[355] = 10'b1111101010;
    16'b0001000010000100: out_v[355] = 10'b0111110101;
    16'b0000000010000000: out_v[355] = 10'b1110110001;
    16'b0101100010000000: out_v[355] = 10'b0100110101;
    16'b0001000010000000: out_v[355] = 10'b1000000111;
    16'b0000000000000000: out_v[355] = 10'b1001010001;
    16'b0100000010000000: out_v[355] = 10'b0011101010;
    16'b0000100010000100: out_v[355] = 10'b0100001011;
    16'b0100100010000100: out_v[355] = 10'b1010000110;
    16'b0101100110000000: out_v[355] = 10'b0100010001;
    16'b0000100000000100: out_v[355] = 10'b0110011010;
    16'b0101100000000000: out_v[355] = 10'b0111111010;
    16'b0101100010000100: out_v[355] = 10'b0110100011;
    16'b0010100010000000: out_v[355] = 10'b0111111001;
    16'b0101000010010000: out_v[355] = 10'b1111000010;
    16'b0000000000000100: out_v[355] = 10'b0110100010;
    16'b0001100010000000: out_v[355] = 10'b0000100110;
    16'b0101100010010000: out_v[355] = 10'b1000010011;
    16'b0010000010000000: out_v[355] = 10'b0001001101;
    16'b0101100110010000: out_v[355] = 10'b1111000011;
    16'b0100000000000000: out_v[355] = 10'b0010101111;
    16'b0101000110000000: out_v[355] = 10'b0011110111;
    16'b0100100000000100: out_v[355] = 10'b0101001001;
    16'b0100000000000100: out_v[355] = 10'b1100111011;
    16'b0100100100000100: out_v[355] = 10'b0001100101;
    16'b0001100000000000: out_v[355] = 10'b1000100101;
    16'b0101100000000100: out_v[355] = 10'b0001101110;
    16'b0001100000000100: out_v[355] = 10'b1011101001;
    16'b0000100100000100: out_v[355] = 10'b1110001011;
    16'b0001000000000100: out_v[355] = 10'b1000010101;
    16'b0100100110000100: out_v[355] = 10'b1100110110;
    16'b0110100010000100: out_v[355] = 10'b0100110100;
    16'b1100100100000100: out_v[355] = 10'b0000101101;
    16'b0001000000000000: out_v[355] = 10'b0101010110;
    16'b0100100100010100: out_v[355] = 10'b0111011011;
    16'b0001000000010100: out_v[355] = 10'b1010100110;
    16'b0101100100000100: out_v[355] = 10'b1110001010;
    16'b0010100010000100: out_v[355] = 10'b1100010110;
    16'b1000100000000100: out_v[355] = 10'b1010101111;
    16'b0100000100000100: out_v[355] = 10'b1010010100;
    16'b0000100100000000: out_v[355] = 10'b0011110110;
    16'b0000101000000100: out_v[355] = 10'b1010011101;
    16'b0110100110000100: out_v[355] = 10'b0110100100;
    16'b0100100100000000: out_v[355] = 10'b1110110111;
    16'b0110100000000100: out_v[355] = 10'b0011110101;
    16'b0001100010000100: out_v[355] = 10'b0001011111;
    16'b0010100000000100: out_v[355] = 10'b1100011001;
    16'b0010100000000000: out_v[355] = 10'b0100100011;
    16'b0110100000000000: out_v[355] = 10'b0100110001;
    16'b0100000100000000: out_v[355] = 10'b0010011110;
    16'b0100000000010000: out_v[355] = 10'b1000011001;
    16'b0101000100000000: out_v[355] = 10'b1001110010;
    16'b0100100000010000: out_v[355] = 10'b1011101011;
    16'b0101000000000000: out_v[355] = 10'b0001011101;
    16'b0110100010000000: out_v[355] = 10'b1110001110;
    16'b0010000000000000: out_v[355] = 10'b1000111100;
    16'b0101100100000000: out_v[355] = 10'b0001101100;
    16'b0000000000010000: out_v[355] = 10'b1010000011;
    16'b0000000010010000: out_v[355] = 10'b1011000001;
    16'b0100000010010000: out_v[355] = 10'b0010011101;
    16'b0100000010000100: out_v[355] = 10'b1100110010;
    16'b0101100100010000: out_v[355] = 10'b0110110010;
    16'b0000001000000100: out_v[355] = 10'b0101101000;
    16'b0101000010000100: out_v[355] = 10'b1011010011;
    16'b0101000000000100: out_v[355] = 10'b0011010110;
    16'b0100001000000100: out_v[355] = 10'b0110010010;
    16'b0101001000000100: out_v[355] = 10'b1110000110;
    16'b0000001000000000: out_v[355] = 10'b1001011010;
    16'b0001001000000100: out_v[355] = 10'b1101011011;
    16'b0000000010010100: out_v[355] = 10'b1101110100;
    16'b0000000000110000: out_v[355] = 10'b1100010111;
    16'b0000000000010100: out_v[355] = 10'b1110001011;
    16'b0000000010110000: out_v[355] = 10'b1111010001;
    16'b0100000000110000: out_v[355] = 10'b0010100011;
    16'b0100100010010100: out_v[355] = 10'b1111110010;
    16'b0100000000010100: out_v[355] = 10'b1000001111;
    16'b0100000010010100: out_v[355] = 10'b0100011111;
    default: out_v[355] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000001000000000: out_v[356] = 10'b1101110010;
    16'b0010000001110000: out_v[356] = 10'b0011111111;
    16'b1001001000010000: out_v[356] = 10'b1111100001;
    16'b0000000000010000: out_v[356] = 10'b1001101010;
    16'b0001000000010000: out_v[356] = 10'b1111100000;
    16'b0011000000110000: out_v[356] = 10'b0110000011;
    16'b0011001000110000: out_v[356] = 10'b1101101100;
    16'b0010000000010000: out_v[356] = 10'b1001110111;
    16'b1011001000000000: out_v[356] = 10'b1110010101;
    16'b0000001000010000: out_v[356] = 10'b0101011111;
    16'b0000000000110000: out_v[356] = 10'b0101101000;
    16'b0011000000010000: out_v[356] = 10'b1101111010;
    16'b0011001000010000: out_v[356] = 10'b0111011010;
    16'b1001001001000000: out_v[356] = 10'b1101000010;
    16'b0000000001010000: out_v[356] = 10'b0000101111;
    16'b1000001000000000: out_v[356] = 10'b1110101110;
    16'b0001001000000000: out_v[356] = 10'b0100010111;
    16'b1001001000000000: out_v[356] = 10'b1100100011;
    16'b1011001000010000: out_v[356] = 10'b0111101010;
    16'b1000001000010000: out_v[356] = 10'b1010101100;
    16'b1001001000110000: out_v[356] = 10'b1010111010;
    16'b0000001000110000: out_v[356] = 10'b1000110110;
    16'b1001000000000000: out_v[356] = 10'b1011010111;
    16'b0010000000110000: out_v[356] = 10'b1110011001;
    16'b0001000000110000: out_v[356] = 10'b0111110000;
    16'b1001001000010001: out_v[356] = 10'b0011000011;
    16'b0001001000010000: out_v[356] = 10'b0010111011;
    16'b1011001000110000: out_v[356] = 10'b1100000011;
    16'b0011000001110000: out_v[356] = 10'b0110101111;
    16'b0000000001000000: out_v[356] = 10'b1000001011;
    16'b1001000000010000: out_v[356] = 10'b1101010010;
    16'b1011001001000000: out_v[356] = 10'b1100110010;
    16'b0000001001000000: out_v[356] = 10'b1010011000;
    16'b1011000000010000: out_v[356] = 10'b0111000100;
    16'b0000000000000000: out_v[356] = 10'b1010100110;
    16'b1001001001010000: out_v[356] = 10'b1011010011;
    16'b0001001000110000: out_v[356] = 10'b1011101100;
    16'b0000000001110000: out_v[356] = 10'b0010101111;
    16'b0000000000100000: out_v[356] = 10'b1001110110;
    16'b1000000000010000: out_v[356] = 10'b0111011100;
    16'b1000000000000000: out_v[356] = 10'b0000110011;
    16'b0000000001100000: out_v[356] = 10'b1100011111;
    16'b1000001000010001: out_v[356] = 10'b1110000100;
    16'b1000000000010001: out_v[356] = 10'b1100110110;
    16'b0000000000000001: out_v[356] = 10'b0100100110;
    16'b1000001000110000: out_v[356] = 10'b1100101001;
    16'b1000001000110010: out_v[356] = 10'b0101100101;
    16'b1000001000000001: out_v[356] = 10'b0011011111;
    16'b1000000000000001: out_v[356] = 10'b0101100111;
    16'b0000000000010001: out_v[356] = 10'b1100110100;
    16'b1000000010010000: out_v[356] = 10'b0010111101;
    16'b1000001010010000: out_v[356] = 10'b1001101110;
    16'b0000001000100000: out_v[356] = 10'b1111000101;
    16'b0000001000010001: out_v[356] = 10'b0010010010;
    16'b1000001000100000: out_v[356] = 10'b1110011101;
    16'b0000000000100010: out_v[356] = 10'b1111101011;
    16'b1000001001010000: out_v[356] = 10'b1001011000;
    16'b1000001000010010: out_v[356] = 10'b0100000110;
    16'b0000001000000001: out_v[356] = 10'b1110100100;
    16'b1000001001000000: out_v[356] = 10'b0111001001;
    16'b0000001000110010: out_v[356] = 10'b1000111101;
    16'b1000000001010000: out_v[356] = 10'b0000111011;
    16'b0000001001010000: out_v[356] = 10'b1101100100;
    16'b1000001010000000: out_v[356] = 10'b1011101011;
    16'b1000000001000000: out_v[356] = 10'b1011110001;
    16'b0000000000010010: out_v[356] = 10'b0101001101;
    16'b1000001011000000: out_v[356] = 10'b1111101011;
    16'b1000000010000000: out_v[356] = 10'b1101001110;
    16'b1000001001100000: out_v[356] = 10'b0011111100;
    16'b1000001001110000: out_v[356] = 10'b1110000100;
    16'b0000000000110010: out_v[356] = 10'b1010011010;
    16'b0001000000000000: out_v[356] = 10'b1010100110;
    16'b1000000000110000: out_v[356] = 10'b1011100100;
    16'b1001000000100000: out_v[356] = 10'b0111101011;
    16'b0000000010000000: out_v[356] = 10'b0010110100;
    16'b0001000000100000: out_v[356] = 10'b0010011000;
    16'b0001000001010000: out_v[356] = 10'b1011001011;
    16'b1001000000110000: out_v[356] = 10'b1010010101;
    16'b0001000010000000: out_v[356] = 10'b1101111111;
    16'b1001001001100000: out_v[356] = 10'b1111100100;
    16'b0001000001000000: out_v[356] = 10'b0100100000;
    16'b0001000001100000: out_v[356] = 10'b0101110000;
    16'b1000000001100000: out_v[356] = 10'b1111100010;
    16'b0001000001110000: out_v[356] = 10'b0111010010;
    16'b0010000000000000: out_v[356] = 10'b1110001011;
    16'b0000001001110000: out_v[356] = 10'b0011111110;
    16'b0010000001010000: out_v[356] = 10'b1011100100;
    16'b1001001000100000: out_v[356] = 10'b0101100111;
    16'b1001000001100000: out_v[356] = 10'b1100110100;
    16'b1001000001000000: out_v[356] = 10'b0011110100;
    16'b1000000000100000: out_v[356] = 10'b1000110101;
    16'b1001000000010001: out_v[356] = 10'b0011110001;
    16'b0011000001010000: out_v[356] = 10'b1001011011;
    16'b0000010000010000: out_v[356] = 10'b0010001010;
    16'b0000000010010000: out_v[356] = 10'b1001100011;
    16'b0000010010010000: out_v[356] = 10'b0010000010;
    16'b0000010000000000: out_v[356] = 10'b1010011001;
    16'b0000010001010000: out_v[356] = 10'b1101001111;
    16'b1010001001010000: out_v[356] = 10'b1000011100;
    default: out_v[356] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0110000000000010: out_v[357] = 10'b0000100100;
    16'b1101000000000010: out_v[357] = 10'b1100001111;
    16'b1111000000000010: out_v[357] = 10'b1101001111;
    16'b1100000000000010: out_v[357] = 10'b0101010110;
    16'b0010000000000000: out_v[357] = 10'b0000011110;
    16'b1001000000000010: out_v[357] = 10'b0101010111;
    16'b1000000000000000: out_v[357] = 10'b0111100111;
    16'b0101000000000010: out_v[357] = 10'b1011001001;
    16'b0000000000000000: out_v[357] = 10'b1011101000;
    16'b1000000000000010: out_v[357] = 10'b0000010001;
    16'b1010000000000010: out_v[357] = 10'b0101010111;
    16'b0001000000000000: out_v[357] = 10'b0010110010;
    16'b1011000000000010: out_v[357] = 10'b1000110011;
    16'b0111000000000010: out_v[357] = 10'b1011001100;
    16'b1010000000000000: out_v[357] = 10'b1001001000;
    16'b0100000000000010: out_v[357] = 10'b0011101000;
    16'b0000000000000010: out_v[357] = 10'b1011011011;
    16'b1110000000000010: out_v[357] = 10'b0001101111;
    16'b1101000000000000: out_v[357] = 10'b1001010011;
    16'b0010000000000010: out_v[357] = 10'b0100000111;
    16'b0011000000000010: out_v[357] = 10'b1100111001;
    16'b1001000000000000: out_v[357] = 10'b0000010110;
    16'b0100000000000000: out_v[357] = 10'b0100010100;
    16'b0101000000000000: out_v[357] = 10'b0010010111;
    16'b0010000010000000: out_v[357] = 10'b0111000100;
    16'b0111000000000000: out_v[357] = 10'b0110010111;
    16'b0110000010000010: out_v[357] = 10'b0100111110;
    16'b1111000001000010: out_v[357] = 10'b1011110011;
    16'b0000000010000010: out_v[357] = 10'b1010001001;
    16'b0010000010000010: out_v[357] = 10'b1110001011;
    16'b0110000000000000: out_v[357] = 10'b0101111100;
    16'b1101000001000010: out_v[357] = 10'b1011110110;
    16'b0000000010000000: out_v[357] = 10'b1010001100;
    16'b0101000001000010: out_v[357] = 10'b0000001110;
    16'b1100000000000000: out_v[357] = 10'b0101010100;
    16'b1001000000100000: out_v[357] = 10'b0001111110;
    16'b1111000000000000: out_v[357] = 10'b0000011011;
    16'b1110000000000000: out_v[357] = 10'b0001011010;
    16'b1011000000000000: out_v[357] = 10'b0111110010;
    16'b1000000000100000: out_v[357] = 10'b0100010010;
    16'b0001000000100000: out_v[357] = 10'b0000101000;
    16'b0001000000000010: out_v[357] = 10'b1100101111;
    16'b1101000000100010: out_v[357] = 10'b1001100011;
    16'b0101000000100010: out_v[357] = 10'b1011101010;
    16'b0000000000100000: out_v[357] = 10'b1100010111;
    16'b1010000010000000: out_v[357] = 10'b0101000101;
    16'b1000000010000000: out_v[357] = 10'b1001100100;
    16'b0100000000100010: out_v[357] = 10'b1111001011;
    16'b0011000000000000: out_v[357] = 10'b0011110100;
    default: out_v[357] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000000000000: out_v[358] = 10'b0010111011;
    16'b0000000000000001: out_v[358] = 10'b0110011011;
    16'b0000010100100001: out_v[358] = 10'b1010000001;
    16'b0000000100100001: out_v[358] = 10'b0001000001;
    16'b0000010100000001: out_v[358] = 10'b0101100011;
    16'b0000000000100000: out_v[358] = 10'b0100110010;
    16'b0000000000100001: out_v[358] = 10'b0001001111;
    16'b0000000100100000: out_v[358] = 10'b1001100000;
    16'b0000010100100000: out_v[358] = 10'b0010011011;
    16'b0000010110100001: out_v[358] = 10'b1001110001;
    16'b0000000100000001: out_v[358] = 10'b1111100011;
    16'b0000010110100000: out_v[358] = 10'b1111110011;
    16'b0000000100000000: out_v[358] = 10'b1010010110;
    16'b0000000010000000: out_v[358] = 10'b0010000111;
    16'b0000000110100000: out_v[358] = 10'b0000011110;
    16'b0000000010100000: out_v[358] = 10'b0100011110;
    16'b0000100000100000: out_v[358] = 10'b1100110101;
    16'b0000000000100010: out_v[358] = 10'b1010111100;
    16'b0000000000101000: out_v[358] = 10'b0000101111;
    16'b0000000000001000: out_v[358] = 10'b1000101100;
    16'b0000010100000000: out_v[358] = 10'b0100111100;
    16'b0000010000000000: out_v[358] = 10'b1010011111;
    16'b0000010010100000: out_v[358] = 10'b1100110110;
    16'b0000010000100000: out_v[358] = 10'b1000101111;
    16'b0000010010000000: out_v[358] = 10'b0010110001;
    16'b0000100100100000: out_v[358] = 10'b1101101010;
    16'b0000100000000000: out_v[358] = 10'b1001000110;
    16'b0000100100100001: out_v[358] = 10'b0101111010;
    16'b0000000010001000: out_v[358] = 10'b1011001111;
    16'b0000010010001000: out_v[358] = 10'b1001001111;
    16'b0000010010000001: out_v[358] = 10'b1110000101;
    16'b0000010011001000: out_v[358] = 10'b1100111110;
    16'b0000010010101000: out_v[358] = 10'b0010110111;
    16'b0000010000101000: out_v[358] = 10'b0110110101;
    16'b0000010000001000: out_v[358] = 10'b1001011110;
    default: out_v[358] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000001000000: out_v[359] = 10'b0100011101;
    16'b0000000000101000: out_v[359] = 10'b0000011110;
    16'b0000000001001001: out_v[359] = 10'b1001010000;
    16'b0000000001001000: out_v[359] = 10'b0100100010;
    16'b0000000001101001: out_v[359] = 10'b0110100111;
    16'b0000000001101000: out_v[359] = 10'b0010101101;
    16'b0000000000000001: out_v[359] = 10'b1100000111;
    16'b0000000000101001: out_v[359] = 10'b0100011101;
    16'b0000100000001001: out_v[359] = 10'b0010111011;
    16'b0000000001100000: out_v[359] = 10'b0110001000;
    16'b0000000000001000: out_v[359] = 10'b0010100110;
    16'b0000000001101010: out_v[359] = 10'b1110000011;
    16'b0000000000001001: out_v[359] = 10'b1101010010;
    16'b0000000001111001: out_v[359] = 10'b1010100111;
    16'b0000100001101001: out_v[359] = 10'b1001001010;
    16'b0000000000100000: out_v[359] = 10'b0100011011;
    16'b0000000001000001: out_v[359] = 10'b1011101000;
    16'b0000000000100001: out_v[359] = 10'b0111010100;
    16'b0000100001001001: out_v[359] = 10'b0101000000;
    16'b0000000000000000: out_v[359] = 10'b1101110000;
    16'b0000000000111001: out_v[359] = 10'b0100001011;
    16'b0000000001100001: out_v[359] = 10'b1010000010;
    16'b0000100001101000: out_v[359] = 10'b0000011100;
    16'b0000110001101001: out_v[359] = 10'b0111011011;
    16'b0000000000101010: out_v[359] = 10'b1001100000;
    16'b0000100000101001: out_v[359] = 10'b1011010010;
    16'b0000100000000000: out_v[359] = 10'b1010001110;
    16'b0000000010000000: out_v[359] = 10'b1011101011;
    16'b0000110000100000: out_v[359] = 10'b0000101100;
    16'b0000100000101000: out_v[359] = 10'b1000011110;
    16'b0000100001001000: out_v[359] = 10'b0000101110;
    16'b0000100000100000: out_v[359] = 10'b0111001100;
    16'b0000010001001000: out_v[359] = 10'b0101101110;
    16'b0000100001100000: out_v[359] = 10'b1010100101;
    16'b0000110000101000: out_v[359] = 10'b0011100111;
    16'b0000100000001000: out_v[359] = 10'b1110100110;
    16'b0000100001000000: out_v[359] = 10'b0101101011;
    16'b0000110001001000: out_v[359] = 10'b1011111111;
    16'b0000110001101000: out_v[359] = 10'b0101010110;
    16'b0000110010100000: out_v[359] = 10'b0100111111;
    16'b0000000010100000: out_v[359] = 10'b0111110100;
    16'b0000010010100000: out_v[359] = 10'b0001111101;
    16'b0000100010100000: out_v[359] = 10'b0011011011;
    16'b0000000011000001: out_v[359] = 10'b1010010100;
    16'b0000010000100001: out_v[359] = 10'b1110011000;
    16'b0000000010100001: out_v[359] = 10'b0111110111;
    16'b0000000001000010: out_v[359] = 10'b0101010101;
    16'b0000010001100001: out_v[359] = 10'b1011000010;
    16'b0000000001000011: out_v[359] = 10'b0001110111;
    16'b0000110001000001: out_v[359] = 10'b0100110010;
    16'b0000100001000001: out_v[359] = 10'b1100101100;
    16'b0000010001000001: out_v[359] = 10'b1010001100;
    16'b0000100011000001: out_v[359] = 10'b0110111111;
    16'b0000000011100000: out_v[359] = 10'b1001010100;
    16'b0000000011000000: out_v[359] = 10'b1100011001;
    16'b0000000011100001: out_v[359] = 10'b1000010111;
    16'b0000000001010001: out_v[359] = 10'b0010011010;
    16'b0000000000100010: out_v[359] = 10'b0000100001;
    16'b0000000000000010: out_v[359] = 10'b0111100100;
    16'b0000100000000001: out_v[359] = 10'b0010110011;
    16'b0000000000001010: out_v[359] = 10'b1110001011;
    16'b0000000000100011: out_v[359] = 10'b1001100111;
    16'b0000000000101011: out_v[359] = 10'b1010100110;
    16'b0000000000000011: out_v[359] = 10'b1000011101;
    16'b0000000100001000: out_v[359] = 10'b1011000000;
    16'b0000000101001000: out_v[359] = 10'b0001110011;
    16'b0000000100101000: out_v[359] = 10'b0111010011;
    16'b0000000100000000: out_v[359] = 10'b0110110010;
    16'b0000000101101000: out_v[359] = 10'b0101001101;
    16'b0000000001110001: out_v[359] = 10'b1110000011;
    16'b0000000001100011: out_v[359] = 10'b1111001011;
    16'b0000010010100001: out_v[359] = 10'b1110100011;
    16'b0000000001001010: out_v[359] = 10'b1110110010;
    16'b0000000001001011: out_v[359] = 10'b0101010011;
    16'b0001010001100001: out_v[359] = 10'b1111001000;
    16'b0000010011100001: out_v[359] = 10'b0010011011;
    default: out_v[359] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100100010000000: out_v[360] = 10'b0001011001;
    16'b0100100010100000: out_v[360] = 10'b0110001001;
    16'b0000101010100000: out_v[360] = 10'b0100000111;
    16'b0000100010010000: out_v[360] = 10'b1001001111;
    16'b0000001010100000: out_v[360] = 10'b0100010100;
    16'b0000100000000000: out_v[360] = 10'b1000111000;
    16'b0000000010000000: out_v[360] = 10'b0100111110;
    16'b0000100010100000: out_v[360] = 10'b0111001011;
    16'b0000001010000000: out_v[360] = 10'b1001010011;
    16'b0000100010101000: out_v[360] = 10'b1010110011;
    16'b0100100010100001: out_v[360] = 10'b0111110101;
    16'b0100100010010000: out_v[360] = 10'b0111110100;
    16'b0101000110100001: out_v[360] = 10'b0011010101;
    16'b0100000010100001: out_v[360] = 10'b1010111111;
    16'b0000100010000000: out_v[360] = 10'b0011100011;
    16'b0100000010101001: out_v[360] = 10'b0111100010;
    16'b0000100010101001: out_v[360] = 10'b0101100001;
    16'b0101001110100001: out_v[360] = 10'b0101001011;
    16'b0100001010100000: out_v[360] = 10'b1111011111;
    16'b0000100011100000: out_v[360] = 10'b0100110001;
    16'b0000100010001000: out_v[360] = 10'b0010111111;
    16'b0100100010101000: out_v[360] = 10'b1010101110;
    16'b0000100000100000: out_v[360] = 10'b1011011001;
    16'b0000100010100001: out_v[360] = 10'b0101111011;
    16'b0000101010000000: out_v[360] = 10'b0001010001;
    16'b0100101010100000: out_v[360] = 10'b0010111111;
    16'b0100000010000000: out_v[360] = 10'b1100100101;
    16'b0000000010101001: out_v[360] = 10'b1011011110;
    16'b0000100011000000: out_v[360] = 10'b1111000001;
    16'b0101100110100001: out_v[360] = 10'b1011111011;
    16'b0100100010101001: out_v[360] = 10'b0101010110;
    16'b0000100010011000: out_v[360] = 10'b1011001111;
    16'b0100000110100001: out_v[360] = 10'b0101110110;
    16'b0100001010100001: out_v[360] = 10'b0011011110;
    16'b0100000010100000: out_v[360] = 10'b0110011111;
    16'b0100100010000001: out_v[360] = 10'b0011111100;
    16'b0100100010001000: out_v[360] = 10'b0111100110;
    16'b0000100010110000: out_v[360] = 10'b1111010010;
    16'b0000000011010000: out_v[360] = 10'b1100110010;
    16'b0000000010010000: out_v[360] = 10'b0100101110;
    16'b0100000000000000: out_v[360] = 10'b0111110001;
    16'b0100000000000001: out_v[360] = 10'b0101011011;
    16'b0100000000001000: out_v[360] = 10'b1010001111;
    16'b0000000000000000: out_v[360] = 10'b1111101110;
    16'b0000000000001000: out_v[360] = 10'b0011000110;
    16'b0000000000000001: out_v[360] = 10'b0110110101;
    16'b0000000011000000: out_v[360] = 10'b1010110010;
    16'b0000000010010100: out_v[360] = 10'b0011110101;
    16'b0100100000000000: out_v[360] = 10'b1111100110;
    16'b0000000010001000: out_v[360] = 10'b1010001010;
    16'b0000000000010000: out_v[360] = 10'b1010000110;
    16'b0000100000000001: out_v[360] = 10'b0011101010;
    16'b0100000000010000: out_v[360] = 10'b1101010111;
    16'b0100100000000001: out_v[360] = 10'b0110111111;
    16'b0001000100010001: out_v[360] = 10'b1010001111;
    16'b0000000110010001: out_v[360] = 10'b0001011000;
    16'b0000000010011001: out_v[360] = 10'b1111010001;
    16'b0001000110010001: out_v[360] = 10'b1100110101;
    16'b0001000110011001: out_v[360] = 10'b0110100011;
    16'b0001000110001001: out_v[360] = 10'b0100011111;
    16'b0000000010011000: out_v[360] = 10'b1100100010;
    16'b0101000100010001: out_v[360] = 10'b0100110111;
    16'b0000000000001001: out_v[360] = 10'b1001100110;
    16'b0000000110011001: out_v[360] = 10'b1111111011;
    16'b0001000110101001: out_v[360] = 10'b0001011100;
    16'b0000000000010001: out_v[360] = 10'b1110011000;
    16'b0000000000011001: out_v[360] = 10'b1111000100;
    16'b0000000010001001: out_v[360] = 10'b1110010100;
    16'b0101000110010001: out_v[360] = 10'b1001011100;
    16'b0101000110011001: out_v[360] = 10'b1111110011;
    16'b0001000110000001: out_v[360] = 10'b1010100101;
    16'b0000000000011000: out_v[360] = 10'b1000110101;
    16'b0000000010010001: out_v[360] = 10'b1101001101;
    16'b0000000010000001: out_v[360] = 10'b1001111100;
    16'b0000000110001001: out_v[360] = 10'b1010110010;
    16'b0000000010100000: out_v[360] = 10'b1100011110;
    16'b0001000100000001: out_v[360] = 10'b1100100100;
    16'b0001000100000000: out_v[360] = 10'b1001101100;
    16'b0100100000010001: out_v[360] = 10'b0010111011;
    16'b0101100100000001: out_v[360] = 10'b1010001000;
    16'b0000100110011001: out_v[360] = 10'b1111110101;
    16'b0101100100010001: out_v[360] = 10'b1111001011;
    16'b0101100110000001: out_v[360] = 10'b0000100010;
    16'b0101000100000001: out_v[360] = 10'b1001011001;
    16'b0000100010011001: out_v[360] = 10'b0111010110;
    16'b0101100110010001: out_v[360] = 10'b0011001000;
    16'b0101100100000000: out_v[360] = 10'b1100110011;
    16'b0001100110010001: out_v[360] = 10'b1011101101;
    16'b0100100000010000: out_v[360] = 10'b1111000111;
    16'b0000100010000001: out_v[360] = 10'b0111100011;
    16'b0100000010010000: out_v[360] = 10'b0001001001;
    16'b0101100100010000: out_v[360] = 10'b0101101011;
    16'b0100100110010001: out_v[360] = 10'b1000001011;
    16'b0101100110011001: out_v[360] = 10'b1111001000;
    16'b0100000010010001: out_v[360] = 10'b0111110010;
    16'b0000100010010001: out_v[360] = 10'b1000011101;
    16'b0000100000010000: out_v[360] = 10'b1010000100;
    16'b0100100010010001: out_v[360] = 10'b1011000010;
    16'b0100100010011001: out_v[360] = 10'b1110011010;
    16'b0100000110010001: out_v[360] = 10'b1001001011;
    16'b0101000110000001: out_v[360] = 10'b0001101110;
    16'b0001100110011001: out_v[360] = 10'b0100110011;
    16'b0000100010001001: out_v[360] = 10'b1010001110;
    16'b0101000100010000: out_v[360] = 10'b0011000011;
    16'b0100100110011001: out_v[360] = 10'b1110110110;
    16'b0101100110001001: out_v[360] = 10'b1001110001;
    16'b0101100110110001: out_v[360] = 10'b0111111110;
    16'b0001000100010000: out_v[360] = 10'b0110010010;
    16'b0000001000000000: out_v[360] = 10'b0100111011;
    16'b0000100000010001: out_v[360] = 10'b0101011001;
    16'b0000000100010000: out_v[360] = 10'b0010010000;
    16'b0000101000010000: out_v[360] = 10'b0101011110;
    16'b0000001000010000: out_v[360] = 10'b0011110101;
    16'b0000100000110000: out_v[360] = 10'b0001111000;
    16'b0001000100110000: out_v[360] = 10'b1111111001;
    16'b0000100100010000: out_v[360] = 10'b0000110011;
    16'b0001100100010000: out_v[360] = 10'b0110111010;
    16'b0000000001010000: out_v[360] = 10'b1101010010;
    16'b0000000000110000: out_v[360] = 10'b1010100111;
    16'b0000001000110000: out_v[360] = 10'b1000011011;
    16'b0000100001010000: out_v[360] = 10'b1100111000;
    16'b0100100000110000: out_v[360] = 10'b0011110101;
    16'b0100101000010000: out_v[360] = 10'b0001011001;
    16'b0100100100010000: out_v[360] = 10'b1101110111;
    16'b0000100011010000: out_v[360] = 10'b0101000010;
    16'b0100100011000000: out_v[360] = 10'b1011011100;
    16'b0100100011010000: out_v[360] = 10'b0010111111;
    16'b0101100110010000: out_v[360] = 10'b1111100101;
    16'b0000100000011001: out_v[360] = 10'b1011001101;
    16'b0000100000111001: out_v[360] = 10'b1010101111;
    16'b0000100000001000: out_v[360] = 10'b1111010001;
    16'b0000100000001001: out_v[360] = 10'b1110001111;
    16'b0000100010111001: out_v[360] = 10'b1110110110;
    16'b0000100000011000: out_v[360] = 10'b1110101010;
    16'b0000100000110001: out_v[360] = 10'b0000001110;
    16'b0000000000111001: out_v[360] = 10'b1101011110;
    16'b0000100010111000: out_v[360] = 10'b1001101110;
    16'b0000100000111000: out_v[360] = 10'b1110000001;
    16'b0000100011110000: out_v[360] = 10'b0011000010;
    16'b0000000000110001: out_v[360] = 10'b1010101111;
    16'b0000100001000000: out_v[360] = 10'b1110011111;
    16'b0000000010111001: out_v[360] = 10'b1101011011;
    16'b0001000100110001: out_v[360] = 10'b0101101000;
    16'b0100100000100000: out_v[360] = 10'b1000010100;
    16'b0100000100010000: out_v[360] = 10'b1010100011;
    16'b0000000000100000: out_v[360] = 10'b1011000110;
    16'b0000100010010100: out_v[360] = 10'b1011000110;
    16'b0100000000100000: out_v[360] = 10'b1011010110;
    16'b0100100010011000: out_v[360] = 10'b0100010101;
    16'b0100100100010001: out_v[360] = 10'b1110001011;
    16'b0001100100000001: out_v[360] = 10'b1110000001;
    16'b0100000000010001: out_v[360] = 10'b0111011011;
    16'b0100100010001001: out_v[360] = 10'b1111010101;
    16'b0100100100000001: out_v[360] = 10'b1011010101;
    16'b0100100000001001: out_v[360] = 10'b1010100111;
    16'b0000100000010100: out_v[360] = 10'b0101110110;
    16'b0100000000110000: out_v[360] = 10'b1010110011;
    default: out_v[360] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100110000010000: out_v[361] = 10'b0111000010;
    16'b0100100010000000: out_v[361] = 10'b1010100011;
    16'b0100000010000000: out_v[361] = 10'b1110110001;
    16'b0100110000000000: out_v[361] = 10'b0011100011;
    16'b0000000011000000: out_v[361] = 10'b1100011101;
    16'b0100100000000000: out_v[361] = 10'b1010000111;
    16'b0000000010000000: out_v[361] = 10'b0110110001;
    16'b0100000011010000: out_v[361] = 10'b0000010101;
    16'b0101110100000000: out_v[361] = 10'b1100101101;
    16'b0000100010000000: out_v[361] = 10'b1111001110;
    16'b0101100000000000: out_v[361] = 10'b1000000110;
    16'b0100000010010000: out_v[361] = 10'b0110100111;
    16'b0100100000010000: out_v[361] = 10'b0001111101;
    16'b0000100000000000: out_v[361] = 10'b0010101111;
    16'b0100000011000000: out_v[361] = 10'b1011011010;
    16'b0100100010010000: out_v[361] = 10'b0001110011;
    16'b0100100011010000: out_v[361] = 10'b1110000000;
    16'b0100000000010000: out_v[361] = 10'b0010011001;
    16'b0110100010000000: out_v[361] = 10'b0011001001;
    16'b0000000010010000: out_v[361] = 10'b1010100100;
    16'b0100100011000000: out_v[361] = 10'b1111111011;
    16'b0100110110000000: out_v[361] = 10'b1100011010;
    16'b0100000000000000: out_v[361] = 10'b1001111001;
    16'b0101110000000000: out_v[361] = 10'b0111000011;
    16'b0100110010000000: out_v[361] = 10'b1010011011;
    16'b0100110010010000: out_v[361] = 10'b1110011111;
    16'b0100110100000000: out_v[361] = 10'b1110111000;
    16'b0101100010000000: out_v[361] = 10'b1011110100;
    16'b0101010100000000: out_v[361] = 10'b0010101010;
    16'b0000000000000000: out_v[361] = 10'b0011101011;
    16'b0000000100000000: out_v[361] = 10'b0001001111;
    16'b0000000100010000: out_v[361] = 10'b1101000101;
    16'b0100000100000000: out_v[361] = 10'b0101000101;
    16'b0100010100000000: out_v[361] = 10'b1010000110;
    16'b0000000000010000: out_v[361] = 10'b1011000010;
    16'b0000010100000000: out_v[361] = 10'b1011000100;
    16'b0001010100000000: out_v[361] = 10'b1100000110;
    16'b0000000000001000: out_v[361] = 10'b0010010011;
    16'b0101000100000000: out_v[361] = 10'b1110010100;
    16'b0101010100010000: out_v[361] = 10'b1001100110;
    16'b0101010100001000: out_v[361] = 10'b1110100001;
    16'b0101100000001000: out_v[361] = 10'b1110001111;
    16'b0001011100001000: out_v[361] = 10'b1011001001;
    16'b0101011100001000: out_v[361] = 10'b0111111101;
    16'b0001010100001000: out_v[361] = 10'b0001011011;
    16'b0100010110000000: out_v[361] = 10'b1001000110;
    16'b0101000000000000: out_v[361] = 10'b1000011000;
    16'b0101011100000000: out_v[361] = 10'b0011110001;
    16'b0001010100010000: out_v[361] = 10'b0100001011;
    16'b0101010110000000: out_v[361] = 10'b1010000111;
    16'b0100010100010000: out_v[361] = 10'b1010000111;
    16'b0100010100001000: out_v[361] = 10'b1000110100;
    16'b0100010101000000: out_v[361] = 10'b1000110011;
    16'b0101010101000000: out_v[361] = 10'b0111001100;
    16'b0101000000010000: out_v[361] = 10'b0000011001;
    16'b0101010100000001: out_v[361] = 10'b1001110101;
    16'b0001011100000000: out_v[361] = 10'b1110111101;
    16'b0101000000001000: out_v[361] = 10'b0110001010;
    16'b0101110100001000: out_v[361] = 10'b0110111000;
    16'b0000010101000000: out_v[361] = 10'b1011010101;
    16'b0000010100001000: out_v[361] = 10'b0111011100;
    16'b0101000100010000: out_v[361] = 10'b0001111111;
    16'b0001010101000000: out_v[361] = 10'b0101101110;
    16'b0001000000000000: out_v[361] = 10'b1010100110;
    16'b0101100000010000: out_v[361] = 10'b0010111110;
    16'b0001100000000001: out_v[361] = 10'b1011101110;
    16'b0001100000010000: out_v[361] = 10'b1001001101;
    16'b0101110100010000: out_v[361] = 10'b0101011010;
    16'b0001000000010000: out_v[361] = 10'b0001001100;
    16'b0001100000000000: out_v[361] = 10'b0011111100;
    16'b0101100000000001: out_v[361] = 10'b1010011010;
    16'b0000100000010000: out_v[361] = 10'b0000110001;
    16'b0101000000000001: out_v[361] = 10'b0000011011;
    16'b0101100010010000: out_v[361] = 10'b1000100110;
    16'b0000110100000000: out_v[361] = 10'b0011111000;
    16'b0011100000000000: out_v[361] = 10'b1000110101;
    16'b0001100100000000: out_v[361] = 10'b0110011100;
    16'b0001110100000000: out_v[361] = 10'b0001111010;
    16'b0011010100000000: out_v[361] = 10'b1100011011;
    16'b0001110100010000: out_v[361] = 10'b0000010011;
    16'b0101110110000000: out_v[361] = 10'b0001011010;
    16'b0011100100000000: out_v[361] = 10'b0010010011;
    16'b0000010100010000: out_v[361] = 10'b0110111001;
    16'b0001110110000000: out_v[361] = 10'b1100111011;
    16'b0001010110000000: out_v[361] = 10'b0101100110;
    16'b0000110100010000: out_v[361] = 10'b0101010000;
    16'b0001100010000000: out_v[361] = 10'b0010011001;
    16'b0101110110010000: out_v[361] = 10'b0110110000;
    16'b0101100100000000: out_v[361] = 10'b0010001110;
    16'b0001110000000000: out_v[361] = 10'b1111001011;
    16'b0011110100000000: out_v[361] = 10'b0010011101;
    16'b0110100100000000: out_v[361] = 10'b1011011111;
    16'b0110100000000000: out_v[361] = 10'b0001001011;
    16'b0111100000000000: out_v[361] = 10'b0010110110;
    16'b0010110100000000: out_v[361] = 10'b1001111110;
    16'b0010100000000000: out_v[361] = 10'b1000101110;
    16'b0110110100000000: out_v[361] = 10'b1010101010;
    16'b0110000000000000: out_v[361] = 10'b1001110000;
    16'b0110110100010000: out_v[361] = 10'b1001101011;
    16'b0111100000010000: out_v[361] = 10'b1010110100;
    16'b0110100000010000: out_v[361] = 10'b1011011011;
    16'b0100110100010000: out_v[361] = 10'b1101011001;
    16'b0000100100000000: out_v[361] = 10'b0101101010;
    16'b0100100100010000: out_v[361] = 10'b0111001001;
    16'b0100100100000000: out_v[361] = 10'b1001011001;
    16'b0000111100000000: out_v[361] = 10'b1010011111;
    16'b0101111100000000: out_v[361] = 10'b0010101111;
    16'b0001010111000000: out_v[361] = 10'b1001100111;
    16'b0001110000001000: out_v[361] = 10'b1011000110;
    16'b0001110110001000: out_v[361] = 10'b0100111011;
    16'b0100101000000000: out_v[361] = 10'b0101010111;
    16'b0000110100001000: out_v[361] = 10'b1011011001;
    16'b0001110100001000: out_v[361] = 10'b1001000010;
    16'b0100111100000000: out_v[361] = 10'b0101011111;
    16'b0101111000000000: out_v[361] = 10'b1111000110;
    16'b0001110111001000: out_v[361] = 10'b1101100100;
    16'b0100011100000000: out_v[361] = 10'b1011010001;
    16'b0001110111000000: out_v[361] = 10'b1111111011;
    16'b0000011100000000: out_v[361] = 10'b1010111001;
    16'b0001111100000000: out_v[361] = 10'b1110101111;
    16'b0101111110000000: out_v[361] = 10'b0101100010;
    16'b0001111000000000: out_v[361] = 10'b1111001111;
    16'b0001010111001000: out_v[361] = 10'b1011001111;
    16'b0001100010001000: out_v[361] = 10'b1011100100;
    16'b0001111110000000: out_v[361] = 10'b1011111010;
    16'b0101101000000000: out_v[361] = 10'b1111110111;
    16'b0000110110000000: out_v[361] = 10'b0101000011;
    16'b0001110010001000: out_v[361] = 10'b1111001011;
    16'b0001000010000000: out_v[361] = 10'b0111100010;
    16'b0001100000001000: out_v[361] = 10'b1000100111;
    16'b0001000010001000: out_v[361] = 10'b0101000010;
    16'b0000110000001000: out_v[361] = 10'b1101010110;
    16'b0001010110001000: out_v[361] = 10'b1111001011;
    16'b0001000100000000: out_v[361] = 10'b0100000111;
    16'b0111110100010000: out_v[361] = 10'b1100011111;
    16'b0111110100000000: out_v[361] = 10'b0101100110;
    16'b0101100100010000: out_v[361] = 10'b0110100001;
    16'b0111010100000000: out_v[361] = 10'b1111001011;
    16'b0101110000010000: out_v[361] = 10'b1110010010;
    16'b0101010000000000: out_v[361] = 10'b0100110111;
    16'b0101010000010000: out_v[361] = 10'b1100001110;
    default: out_v[361] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1000010001000000: out_v[362] = 10'b1101001001;
    16'b1000000000100000: out_v[362] = 10'b0000111011;
    16'b1000001001100000: out_v[362] = 10'b1101010100;
    16'b1000000001100000: out_v[362] = 10'b1101110010;
    16'b1000010000000000: out_v[362] = 10'b0100010011;
    16'b0000000001000000: out_v[362] = 10'b0100011011;
    16'b0000001001100000: out_v[362] = 10'b0110011001;
    16'b0000001000000000: out_v[362] = 10'b1001100011;
    16'b0000000000100000: out_v[362] = 10'b0101111000;
    16'b0000010001000000: out_v[362] = 10'b0101110111;
    16'b0000000001100000: out_v[362] = 10'b0100101100;
    16'b1000000000000000: out_v[362] = 10'b1010101110;
    16'b0000010000000000: out_v[362] = 10'b0101010101;
    16'b0000000101000000: out_v[362] = 10'b0110100011;
    16'b0000001001000000: out_v[362] = 10'b0001011011;
    16'b0000000000000000: out_v[362] = 10'b1000111011;
    16'b1000010000100000: out_v[362] = 10'b0000011101;
    16'b1000000001000000: out_v[362] = 10'b1010111000;
    16'b1000001000100000: out_v[362] = 10'b1001001011;
    16'b0000011001000000: out_v[362] = 10'b1011101110;
    16'b1000011000100000: out_v[362] = 10'b1110100011;
    16'b1000010000000100: out_v[362] = 10'b0001011111;
    16'b1000010000100100: out_v[362] = 10'b1010000010;
    16'b0000001000100000: out_v[362] = 10'b1000011011;
    16'b1000010001100000: out_v[362] = 10'b0101000100;
    16'b1000000000100100: out_v[362] = 10'b1100110001;
    16'b0000010001100000: out_v[362] = 10'b1001100111;
    16'b1000010001000100: out_v[362] = 10'b1011010100;
    16'b0000011001100000: out_v[362] = 10'b1010101111;
    16'b0000010000000100: out_v[362] = 10'b1100101010;
    16'b0000000000000100: out_v[362] = 10'b1001001011;
    16'b0000100000000110: out_v[362] = 10'b0100001111;
    16'b0000010000100100: out_v[362] = 10'b0111011110;
    16'b0000010000101100: out_v[362] = 10'b1111001110;
    16'b0000010001000100: out_v[362] = 10'b0001010101;
    16'b1000000100000000: out_v[362] = 10'b1100101001;
    16'b0000010001100100: out_v[362] = 10'b1110000101;
    16'b1000010100000100: out_v[362] = 10'b0110001101;
    16'b0000010101000100: out_v[362] = 10'b1001101100;
    16'b0000000001000100: out_v[362] = 10'b1001000111;
    16'b1000000101000100: out_v[362] = 10'b0111011011;
    16'b0000010100000100: out_v[362] = 10'b1010111101;
    16'b1000000000000100: out_v[362] = 10'b0110010001;
    16'b1000010001100100: out_v[362] = 10'b1111010110;
    16'b1000000100000100: out_v[362] = 10'b0111001101;
    16'b1000010101000100: out_v[362] = 10'b1001101010;
    16'b1000000001000100: out_v[362] = 10'b1101000000;
    16'b1000000101000000: out_v[362] = 10'b0110110110;
    16'b0000010101000000: out_v[362] = 10'b1000000111;
    16'b0000000101000100: out_v[362] = 10'b1110000010;
    16'b1000000001100100: out_v[362] = 10'b0001101010;
    16'b1000010101100100: out_v[362] = 10'b0101100111;
    16'b1010000000100000: out_v[362] = 10'b0111001010;
    16'b1000100000000010: out_v[362] = 10'b1010001010;
    16'b1000100001000010: out_v[362] = 10'b0010101100;
    16'b1010000001000000: out_v[362] = 10'b1000011001;
    16'b1010000000000000: out_v[362] = 10'b1101011110;
    16'b1000000000101000: out_v[362] = 10'b0110000111;
    16'b0000000000101100: out_v[362] = 10'b0001111000;
    16'b0000100000000010: out_v[362] = 10'b1010110100;
    16'b1000010000101100: out_v[362] = 10'b0110010000;
    16'b1000100000100010: out_v[362] = 10'b1110000111;
    16'b1000000000101100: out_v[362] = 10'b1011010011;
    16'b0000000000100100: out_v[362] = 10'b1010100101;
    16'b1000100000000110: out_v[362] = 10'b1011000110;
    16'b1000100000100110: out_v[362] = 10'b0010110011;
    16'b1000000001101000: out_v[362] = 10'b1110111111;
    16'b0000011000000100: out_v[362] = 10'b0101100111;
    16'b0000010000100000: out_v[362] = 10'b1001110110;
    16'b1000000000001000: out_v[362] = 10'b1100110011;
    16'b0000100000100110: out_v[362] = 10'b0000100111;
    16'b1000000001001000: out_v[362] = 10'b1110101101;
    16'b0000000000101000: out_v[362] = 10'b1010111111;
    16'b0000001000000100: out_v[362] = 10'b0010100010;
    16'b1000100001100010: out_v[362] = 10'b0011100011;
    16'b1000010101000000: out_v[362] = 10'b0111010111;
    16'b1000010100000000: out_v[362] = 10'b0101000100;
    16'b0000011001000100: out_v[362] = 10'b1001011011;
    16'b0000000100000100: out_v[362] = 10'b1001011001;
    16'b0000010100000000: out_v[362] = 10'b1101010100;
    16'b1000110000000110: out_v[362] = 10'b0111110000;
    16'b0000011000100100: out_v[362] = 10'b0011011001;
    16'b0000110000100110: out_v[362] = 10'b1100000011;
    16'b0000110000000110: out_v[362] = 10'b1101000101;
    default: out_v[362] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000000100011: out_v[363] = 10'b1100101011;
    16'b0010001000100011: out_v[363] = 10'b1111111010;
    16'b0010000000100011: out_v[363] = 10'b0101111101;
    16'b0000000001100011: out_v[363] = 10'b0001010111;
    16'b1000000000000011: out_v[363] = 10'b1001100000;
    16'b1000000000100000: out_v[363] = 10'b0010001001;
    16'b0000000000100010: out_v[363] = 10'b1010000010;
    16'b0000000000000001: out_v[363] = 10'b0101010011;
    16'b0000000000100000: out_v[363] = 10'b0011011111;
    16'b0010010000100010: out_v[363] = 10'b1000001011;
    16'b0000001001100011: out_v[363] = 10'b1011111011;
    16'b0000000000100001: out_v[363] = 10'b0101011001;
    16'b1000001001000011: out_v[363] = 10'b0111010000;
    16'b0010010000100011: out_v[363] = 10'b1011000011;
    16'b0010000000000011: out_v[363] = 10'b1000100001;
    16'b0000000000000010: out_v[363] = 10'b0101110100;
    16'b0010000001100010: out_v[363] = 10'b1010001111;
    16'b1000000000100010: out_v[363] = 10'b0011011011;
    16'b1010000001100011: out_v[363] = 10'b1000011111;
    16'b1000000000100011: out_v[363] = 10'b1100111010;
    16'b1000000001100011: out_v[363] = 10'b1110100110;
    16'b0010000000100001: out_v[363] = 10'b1000110011;
    16'b0000000000000011: out_v[363] = 10'b1011000101;
    16'b0010000000100000: out_v[363] = 10'b1001000111;
    16'b0010000000100010: out_v[363] = 10'b0000010101;
    16'b1000001000100010: out_v[363] = 10'b0110101111;
    16'b0010010000000010: out_v[363] = 10'b0001111011;
    16'b1010000000100011: out_v[363] = 10'b1101011011;
    16'b0000001000100011: out_v[363] = 10'b0110000001;
    16'b1000001000100011: out_v[363] = 10'b1110101111;
    16'b1000001001100011: out_v[363] = 10'b1000100001;
    16'b0010010000100000: out_v[363] = 10'b1101110001;
    16'b1000000000000010: out_v[363] = 10'b1011011011;
    16'b0010000001100011: out_v[363] = 10'b0001110111;
    16'b1010000000000011: out_v[363] = 10'b1101000011;
    16'b0010000000000010: out_v[363] = 10'b0000110111;
    16'b1000000000100001: out_v[363] = 10'b0110010100;
    16'b1010010000100011: out_v[363] = 10'b0001111001;
    16'b1010001001100011: out_v[363] = 10'b1111000001;
    16'b1000001001100010: out_v[363] = 10'b0010110011;
    16'b1000001001000010: out_v[363] = 10'b0001010101;
    16'b0010010000100001: out_v[363] = 10'b0110000111;
    16'b1000000001000001: out_v[363] = 10'b1010111000;
    16'b0000001001000000: out_v[363] = 10'b1000100010;
    16'b0000000001000000: out_v[363] = 10'b1101001001;
    16'b0000000000000000: out_v[363] = 10'b0011000011;
    16'b0010001000000000: out_v[363] = 10'b1000101000;
    16'b0000001000000000: out_v[363] = 10'b1000111101;
    16'b0000001000000001: out_v[363] = 10'b0100110001;
    16'b0010001000000001: out_v[363] = 10'b0000011111;
    16'b0010011000000001: out_v[363] = 10'b1000011010;
    16'b1000001001000000: out_v[363] = 10'b0011010011;
    16'b1000001000000001: out_v[363] = 10'b1100000110;
    16'b0000000001000010: out_v[363] = 10'b1011110100;
    16'b1010001000000001: out_v[363] = 10'b1101100110;
    16'b0000001001000010: out_v[363] = 10'b0101001010;
    16'b1010011000000001: out_v[363] = 10'b0101110011;
    16'b0010010001000000: out_v[363] = 10'b0011011101;
    16'b0010011001000001: out_v[363] = 10'b0010111101;
    16'b1010010001000011: out_v[363] = 10'b0011110111;
    16'b1010010000000001: out_v[363] = 10'b1111000110;
    16'b0010010001000001: out_v[363] = 10'b0111011001;
    16'b1000000001100010: out_v[363] = 10'b1100010110;
    16'b1000000001000010: out_v[363] = 10'b0010111100;
    16'b0010010000000000: out_v[363] = 10'b0001110100;
    16'b1010000000000000: out_v[363] = 10'b0110100101;
    16'b1010000000000001: out_v[363] = 10'b0110100111;
    16'b1010010000000011: out_v[363] = 10'b1110000111;
    16'b1010010001000010: out_v[363] = 10'b1000101110;
    16'b0010000001000001: out_v[363] = 10'b1000110001;
    16'b1000000000000000: out_v[363] = 10'b0111101101;
    16'b0010010000000001: out_v[363] = 10'b0010011100;
    16'b0010001001000011: out_v[363] = 10'b1000101110;
    16'b1010000001100010: out_v[363] = 10'b0011110110;
    16'b1010010001100011: out_v[363] = 10'b0110110100;
    16'b1000000001000011: out_v[363] = 10'b1000011000;
    16'b1010010001100010: out_v[363] = 10'b0101101010;
    16'b0010011001000011: out_v[363] = 10'b1001101100;
    16'b0010000000000001: out_v[363] = 10'b1100001010;
    16'b1000010001000010: out_v[363] = 10'b1111110111;
    16'b1010000001000011: out_v[363] = 10'b1011110011;
    16'b1010000001000010: out_v[363] = 10'b0011110111;
    16'b0000000001000011: out_v[363] = 10'b0010111100;
    16'b1010010001000000: out_v[363] = 10'b1010110001;
    16'b1010010001000001: out_v[363] = 10'b1000111011;
    16'b0010010001000011: out_v[363] = 10'b0010110111;
    16'b0010000001000011: out_v[363] = 10'b0000111011;
    16'b1010011001000010: out_v[363] = 10'b1100010000;
    16'b1010000001000000: out_v[363] = 10'b1000101110;
    16'b1010010000100001: out_v[363] = 10'b1101010110;
    16'b0010011001000000: out_v[363] = 10'b1101000100;
    16'b1010010000000000: out_v[363] = 10'b0111011000;
    16'b0010000001000000: out_v[363] = 10'b0001011101;
    16'b0010000000000000: out_v[363] = 10'b0110110100;
    16'b1000000001000000: out_v[363] = 10'b1001000101;
    16'b0010000001000010: out_v[363] = 10'b0111101001;
    16'b0010010001000010: out_v[363] = 10'b1001011010;
    16'b1010011000000000: out_v[363] = 10'b1001001011;
    16'b1000001000100001: out_v[363] = 10'b1100101010;
    16'b1010011001000001: out_v[363] = 10'b0010011011;
    16'b0010011000000000: out_v[363] = 10'b0011111001;
    16'b1010011001000011: out_v[363] = 10'b1110001010;
    16'b1010001000000000: out_v[363] = 10'b1100111001;
    16'b1000011000000001: out_v[363] = 10'b0110011000;
    16'b0010001001000001: out_v[363] = 10'b0000001111;
    16'b1010011001000000: out_v[363] = 10'b0110010101;
    16'b1010001000100001: out_v[363] = 10'b0011110110;
    16'b1010001000000011: out_v[363] = 10'b1000101110;
    16'b1010011000000011: out_v[363] = 10'b1000111000;
    16'b1010011000100001: out_v[363] = 10'b1101101111;
    16'b0010011000000011: out_v[363] = 10'b1010101101;
    16'b1010000001000001: out_v[363] = 10'b1101000110;
    16'b1010001001000000: out_v[363] = 10'b0110010010;
    16'b1010001001000001: out_v[363] = 10'b0101011011;
    16'b1000001000000000: out_v[363] = 10'b1101100100;
    16'b0010011000000010: out_v[363] = 10'b1110101100;
    16'b1000001001000001: out_v[363] = 10'b0011010001;
    16'b1010001001000011: out_v[363] = 10'b0001101010;
    16'b1000000001100000: out_v[363] = 10'b0001111000;
    16'b1000000000000001: out_v[363] = 10'b0110011111;
    16'b1000001000100000: out_v[363] = 10'b1101010100;
    16'b1000000001100001: out_v[363] = 10'b0100011101;
    16'b1010000001100000: out_v[363] = 10'b0110100101;
    16'b1010000001100001: out_v[363] = 10'b1110110010;
    16'b0000001000100000: out_v[363] = 10'b1100100101;
    16'b1000001000000011: out_v[363] = 10'b0010111100;
    16'b0000000001000001: out_v[363] = 10'b0001111101;
    16'b1000001000000010: out_v[363] = 10'b0101101110;
    16'b0000001000100010: out_v[363] = 10'b0010111011;
    16'b0000001001100000: out_v[363] = 10'b0100100010;
    16'b0000001001100010: out_v[363] = 10'b0111000000;
    16'b0000000001100000: out_v[363] = 10'b1000101100;
    16'b0010001000000010: out_v[363] = 10'b0111011100;
    16'b1000000101000011: out_v[363] = 10'b1010111011;
    16'b0010010011000001: out_v[363] = 10'b1111011010;
    16'b0010000011000001: out_v[363] = 10'b0111101001;
    16'b1010010011000011: out_v[363] = 10'b1101110011;
    16'b0010010010000011: out_v[363] = 10'b1010010101;
    16'b1000000100000011: out_v[363] = 10'b1100110111;
    16'b0010010011000011: out_v[363] = 10'b1110111011;
    16'b1010010010000011: out_v[363] = 10'b0101111110;
    16'b0000001001000011: out_v[363] = 10'b0111000011;
    16'b0000000101000011: out_v[363] = 10'b1100111111;
    16'b1000001101000010: out_v[363] = 10'b1111001001;
    16'b1000001101000011: out_v[363] = 10'b1010010111;
    16'b0000001001000001: out_v[363] = 10'b0111000110;
    16'b1000001101000001: out_v[363] = 10'b1111110111;
    16'b0010010000000011: out_v[363] = 10'b0111100001;
    16'b1010000011000001: out_v[363] = 10'b1101100011;
    16'b1010000011000011: out_v[363] = 10'b1110100011;
    16'b0010011001100011: out_v[363] = 10'b0101100010;
    16'b1000100000100000: out_v[363] = 10'b0011110111;
    16'b0000100000000000: out_v[363] = 10'b1011000101;
    16'b1000100000000000: out_v[363] = 10'b0010111011;
    16'b1000100000000001: out_v[363] = 10'b1111111110;
    16'b1000000000010001: out_v[363] = 10'b0110111110;
    16'b1000000000110001: out_v[363] = 10'b0100101011;
    16'b1000100000100001: out_v[363] = 10'b0111111101;
    16'b1010000000100000: out_v[363] = 10'b1011001010;
    16'b1000000000010000: out_v[363] = 10'b0111110111;
    16'b0010001001100001: out_v[363] = 10'b1011110111;
    16'b1010001001100010: out_v[363] = 10'b1100010011;
    16'b0000000001100010: out_v[363] = 10'b1100000010;
    16'b0000000001100001: out_v[363] = 10'b0110100011;
    16'b1000001001100001: out_v[363] = 10'b0001111001;
    16'b0010001001000000: out_v[363] = 10'b0111011000;
    16'b1010011001100000: out_v[363] = 10'b0010000101;
    16'b1010001001100000: out_v[363] = 10'b1001100001;
    16'b1000001001100000: out_v[363] = 10'b1110110010;
    16'b1010011001100011: out_v[363] = 10'b0101000011;
    16'b0010001001100000: out_v[363] = 10'b0111001001;
    16'b1010001001100001: out_v[363] = 10'b0010010101;
    16'b0000001001100001: out_v[363] = 10'b0001110101;
    16'b1010010001100000: out_v[363] = 10'b0111000011;
    16'b1010001001000010: out_v[363] = 10'b0100000011;
    16'b0010000001100001: out_v[363] = 10'b1001110110;
    16'b0010000001100000: out_v[363] = 10'b1100101010;
    16'b1010011001100001: out_v[363] = 10'b0000101111;
    16'b1010011001100010: out_v[363] = 10'b1111010110;
    16'b0010001001100011: out_v[363] = 10'b1111110111;
    16'b0010001001100010: out_v[363] = 10'b1101010110;
    16'b1000100001100000: out_v[363] = 10'b1100100111;
    16'b1000100001000000: out_v[363] = 10'b1101101101;
    16'b1010000000000010: out_v[363] = 10'b1101000110;
    16'b1000101000000000: out_v[363] = 10'b1101000001;
    default: out_v[363] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100000100000000: out_v[364] = 10'b1001001001;
    16'b0100010100100000: out_v[364] = 10'b0100001000;
    16'b0000010100000001: out_v[364] = 10'b0000110101;
    16'b0000010000000010: out_v[364] = 10'b1100100100;
    16'b0000010000000000: out_v[364] = 10'b0100101001;
    16'b0100000100000001: out_v[364] = 10'b0110111010;
    16'b0100000100000010: out_v[364] = 10'b1110101101;
    16'b0100010100000001: out_v[364] = 10'b0100000001;
    16'b0100010000000000: out_v[364] = 10'b0001110111;
    16'b0000000100000001: out_v[364] = 10'b1101111000;
    16'b0100010100000000: out_v[364] = 10'b0100001101;
    16'b0000000100000000: out_v[364] = 10'b1101100011;
    16'b0000010100000000: out_v[364] = 10'b1101001101;
    16'b0100010100100001: out_v[364] = 10'b0000001001;
    16'b0000010100100000: out_v[364] = 10'b1001001111;
    16'b0100000100100000: out_v[364] = 10'b0010101100;
    16'b0100010000000001: out_v[364] = 10'b0101100001;
    16'b0100010100000010: out_v[364] = 10'b1111000101;
    16'b0000010100100010: out_v[364] = 10'b0011010111;
    16'b0000010000000001: out_v[364] = 10'b1100011111;
    16'b0000000000000000: out_v[364] = 10'b1110001110;
    16'b0100000000000000: out_v[364] = 10'b0001110010;
    16'b0000000100100000: out_v[364] = 10'b0011111111;
    16'b0100010000100000: out_v[364] = 10'b0100001111;
    16'b0100010100100010: out_v[364] = 10'b0111000000;
    16'b0100000100100001: out_v[364] = 10'b0100100100;
    16'b0000000000000001: out_v[364] = 10'b1001011001;
    16'b0000000101100010: out_v[364] = 10'b0000010110;
    16'b0000000101000010: out_v[364] = 10'b0010110110;
    16'b0000000000000010: out_v[364] = 10'b0001011001;
    16'b0000000001000010: out_v[364] = 10'b1001001011;
    16'b0100000001000010: out_v[364] = 10'b1011110000;
    16'b0100000101000010: out_v[364] = 10'b0010111110;
    16'b0000000001100010: out_v[364] = 10'b0101011110;
    16'b0000000000100000: out_v[364] = 10'b1111100011;
    16'b0000000001100000: out_v[364] = 10'b1100110111;
    16'b0100000000000010: out_v[364] = 10'b0110011010;
    16'b0100000101100010: out_v[364] = 10'b1100101001;
    16'b0100000101000000: out_v[364] = 10'b1111110101;
    16'b0100000101000011: out_v[364] = 10'b1101110100;
    16'b0100000001100010: out_v[364] = 10'b0101001110;
    16'b0000000001000011: out_v[364] = 10'b0010001001;
    16'b0000010001000010: out_v[364] = 10'b0100100101;
    16'b0100010101100010: out_v[364] = 10'b0101100010;
    16'b0000000101000011: out_v[364] = 10'b0110000100;
    16'b0100000100000011: out_v[364] = 10'b0001001111;
    16'b0100010001100010: out_v[364] = 10'b1010100100;
    16'b0100010101000010: out_v[364] = 10'b0110111100;
    16'b0100010001000010: out_v[364] = 10'b1000100110;
    16'b0100010001000011: out_v[364] = 10'b0011110110;
    16'b0000010001000011: out_v[364] = 10'b0111011100;
    16'b0000010001100010: out_v[364] = 10'b1001111011;
    16'b0100000101001011: out_v[364] = 10'b0110111011;
    16'b0100000101100011: out_v[364] = 10'b1101110110;
    16'b0100010101000011: out_v[364] = 10'b1000110101;
    16'b0100010000100010: out_v[364] = 10'b1110001111;
    16'b0100001101001011: out_v[364] = 10'b1000101111;
    16'b0100010000000010: out_v[364] = 10'b0111100110;
    16'b0100000001000011: out_v[364] = 10'b0001110100;
    16'b0100010001100011: out_v[364] = 10'b1001101101;
    16'b0000000001001011: out_v[364] = 10'b0000001110;
    16'b0100010101100011: out_v[364] = 10'b0011010111;
    16'b0000001001001011: out_v[364] = 10'b1110000101;
    16'b0100000000000001: out_v[364] = 10'b0100100011;
    16'b0100001100001001: out_v[364] = 10'b1100110011;
    16'b0000001100001001: out_v[364] = 10'b1101011011;
    16'b0000001000001001: out_v[364] = 10'b0100000111;
    16'b0010001100001001: out_v[364] = 10'b1011100011;
    16'b0000000100000010: out_v[364] = 10'b1110100000;
    16'b0000000100001001: out_v[364] = 10'b0001011111;
    16'b0110001100001000: out_v[364] = 10'b1100001011;
    16'b0100000100001001: out_v[364] = 10'b0101111010;
    16'b0100000000100000: out_v[364] = 10'b0011101001;
    16'b0100000100100010: out_v[364] = 10'b0100100000;
    16'b0000000000000011: out_v[364] = 10'b0011100001;
    16'b0000000001000111: out_v[364] = 10'b0101101000;
    16'b0100000000000011: out_v[364] = 10'b0101111110;
    16'b0000000000100010: out_v[364] = 10'b0101110010;
    16'b0000010101100010: out_v[364] = 10'b1111011000;
    16'b0000000000100001: out_v[364] = 10'b1011011011;
    16'b0000000000000111: out_v[364] = 10'b1101000101;
    16'b0000000100100010: out_v[364] = 10'b0111100001;
    16'b0000000001100011: out_v[364] = 10'b1001110101;
    16'b0000000000000101: out_v[364] = 10'b0001110110;
    16'b0000000000000100: out_v[364] = 10'b1010010001;
    16'b0000000000100011: out_v[364] = 10'b1011001110;
    16'b0000010101000010: out_v[364] = 10'b1010111010;
    16'b0000010100000010: out_v[364] = 10'b0000010011;
    16'b0000000100100001: out_v[364] = 10'b0100101110;
    16'b0100000001000000: out_v[364] = 10'b0110000101;
    16'b0000010000000011: out_v[364] = 10'b0101001111;
    16'b0000000001000000: out_v[364] = 10'b0111011010;
    16'b0100110001100010: out_v[364] = 10'b1111101101;
    16'b0100100001000010: out_v[364] = 10'b1010101101;
    16'b0000000100000011: out_v[364] = 10'b1000111000;
    16'b0001000000000000: out_v[364] = 10'b0010001001;
    16'b0000001000001101: out_v[364] = 10'b0011000010;
    16'b0001000000000001: out_v[364] = 10'b1001011000;
    16'b0000000000001011: out_v[364] = 10'b0110110011;
    16'b0000001000001011: out_v[364] = 10'b0010110100;
    16'b0000001101001011: out_v[364] = 10'b1111000011;
    16'b0000001100001011: out_v[364] = 10'b0101110000;
    16'b0000000100001011: out_v[364] = 10'b0001010001;
    16'b0000000000001001: out_v[364] = 10'b0111100110;
    16'b0001000000000101: out_v[364] = 10'b1101000011;
    16'b0100000000100010: out_v[364] = 10'b1111000100;
    16'b0100000100000101: out_v[364] = 10'b0110011010;
    16'b0000000001000110: out_v[364] = 10'b1000100101;
    default: out_v[364] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000000000000: out_v[365] = 10'b0111010011;
    16'b0000000100110000: out_v[365] = 10'b0100010101;
    16'b0000000100100000: out_v[365] = 10'b1110100011;
    16'b0000000100100010: out_v[365] = 10'b1100100001;
    16'b0000000000100010: out_v[365] = 10'b1110000101;
    16'b0000000000110000: out_v[365] = 10'b0000010101;
    16'b0000000000100000: out_v[365] = 10'b1010010110;
    16'b0000000000000010: out_v[365] = 10'b0101010011;
    16'b0010000100100000: out_v[365] = 10'b1000110011;
    16'b0000000100000010: out_v[365] = 10'b1000011111;
    16'b0000000100000000: out_v[365] = 10'b1110001111;
    16'b0000000100110010: out_v[365] = 10'b1011011101;
    16'b0000000100010000: out_v[365] = 10'b1110100001;
    16'b0010000100100010: out_v[365] = 10'b0100110001;
    16'b0010000100000000: out_v[365] = 10'b1100111010;
    16'b0010000000100000: out_v[365] = 10'b0101111000;
    16'b0010000100110000: out_v[365] = 10'b0110101010;
    16'b0010000100010000: out_v[365] = 10'b1110110001;
    16'b0010000000000000: out_v[365] = 10'b1101011100;
    16'b0010000000000010: out_v[365] = 10'b0111000100;
    16'b0010000100000010: out_v[365] = 10'b1011001101;
    16'b0010000000110000: out_v[365] = 10'b1101001011;
    16'b0011000000000000: out_v[365] = 10'b1011010100;
    16'b0010000000100010: out_v[365] = 10'b1111001110;
    16'b0001000000000010: out_v[365] = 10'b0110111100;
    16'b0000010000000000: out_v[365] = 10'b1110000010;
    16'b1000000000000010: out_v[365] = 10'b0111011010;
    16'b1010000000000000: out_v[365] = 10'b0010100111;
    16'b0011000000000010: out_v[365] = 10'b1010011001;
    16'b1000000000000000: out_v[365] = 10'b1101110100;
    16'b0000000000110010: out_v[365] = 10'b0001011101;
    16'b1010000000000010: out_v[365] = 10'b1001001011;
    16'b0001000000000000: out_v[365] = 10'b0101100100;
    16'b0000010100000000: out_v[365] = 10'b0100011110;
    16'b0000000000001000: out_v[365] = 10'b1011001010;
    16'b0010000100001000: out_v[365] = 10'b1111011011;
    16'b0010010100000000: out_v[365] = 10'b1101101101;
    16'b0010010000000000: out_v[365] = 10'b1100011000;
    16'b0010010100001000: out_v[365] = 10'b1100100110;
    16'b0010010000001000: out_v[365] = 10'b0001101010;
    16'b0010010100100000: out_v[365] = 10'b1001101010;
    16'b0010000100110010: out_v[365] = 10'b0111011010;
    16'b0010000000001000: out_v[365] = 10'b1001001010;
    16'b0000000000010000: out_v[365] = 10'b0011111010;
    16'b0000010000001000: out_v[365] = 10'b0001110100;
    16'b0000010000100000: out_v[365] = 10'b1010100001;
    16'b0010000000010000: out_v[365] = 10'b0101110010;
    16'b0000000100010010: out_v[365] = 10'b0110110000;
    16'b0010000100010010: out_v[365] = 10'b1000100011;
    16'b0000010100100000: out_v[365] = 10'b0010110100;
    16'b0000010010000000: out_v[365] = 10'b0111001010;
    16'b0000100000000000: out_v[365] = 10'b1101111101;
    16'b0000110000000000: out_v[365] = 10'b1001111001;
    16'b0010010000100000: out_v[365] = 10'b1101011010;
    default: out_v[365] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000100001000: out_v[366] = 10'b0001110110;
    16'b0001010000101011: out_v[366] = 10'b0010100011;
    16'b1001010000101011: out_v[366] = 10'b1011101011;
    16'b0001000001001000: out_v[366] = 10'b0100011111;
    16'b0001010000100010: out_v[366] = 10'b0000111110;
    16'b0001000000100011: out_v[366] = 10'b0010111011;
    16'b0001000000101010: out_v[366] = 10'b1100110111;
    16'b0000000100000000: out_v[366] = 10'b1011000010;
    16'b0001100101001000: out_v[366] = 10'b1001001111;
    16'b0001010000001001: out_v[366] = 10'b1011111101;
    16'b0001010100101011: out_v[366] = 10'b1011010111;
    16'b0001000000001000: out_v[366] = 10'b1000001001;
    16'b0001010000100011: out_v[366] = 10'b0010011011;
    16'b0001000000101011: out_v[366] = 10'b0010011001;
    16'b0001010000101010: out_v[366] = 10'b0110111011;
    16'b1001000111001000: out_v[366] = 10'b0100010101;
    16'b0001000100001000: out_v[366] = 10'b0111010110;
    16'b0000000101001000: out_v[366] = 10'b1001001111;
    16'b1001010100101011: out_v[366] = 10'b1011110101;
    16'b0001010010101011: out_v[366] = 10'b1001011110;
    16'b0000000000100001: out_v[366] = 10'b1010101001;
    16'b0001010001101011: out_v[366] = 10'b1000010011;
    16'b1001000101001000: out_v[366] = 10'b1111100011;
    16'b0001000000101001: out_v[366] = 10'b1111011010;
    16'b0001110001101011: out_v[366] = 10'b1111000010;
    16'b1001100111001000: out_v[366] = 10'b1110000001;
    16'b0001000101001000: out_v[366] = 10'b0100110010;
    16'b0001010101101011: out_v[366] = 10'b1000100111;
    16'b0000000101000000: out_v[366] = 10'b1001100001;
    16'b0001010000101001: out_v[366] = 10'b0110111111;
    16'b0001000000000000: out_v[366] = 10'b0011101010;
    16'b0000010000101011: out_v[366] = 10'b1010110101;
    16'b0001010001100011: out_v[366] = 10'b0101111010;
    16'b0000000000000000: out_v[366] = 10'b0010101100;
    16'b0001000100001001: out_v[366] = 10'b1010110111;
    16'b0001000000100001: out_v[366] = 10'b0011101011;
    16'b1000010000101011: out_v[366] = 10'b1000110111;
    16'b0000000000001000: out_v[366] = 10'b0010110111;
    16'b0000000000100011: out_v[366] = 10'b0110011001;
    16'b0001000000001001: out_v[366] = 10'b1111110011;
    16'b0000100010001000: out_v[366] = 10'b1100110101;
    16'b0000100000001000: out_v[366] = 10'b1101000111;
    16'b0000100001000000: out_v[366] = 10'b0011100011;
    16'b0000100000000000: out_v[366] = 10'b1101000100;
    16'b1000100010001000: out_v[366] = 10'b1101011111;
    16'b0000100101001000: out_v[366] = 10'b0101001011;
    16'b0000100101000000: out_v[366] = 10'b0101111100;
    16'b0000100100001000: out_v[366] = 10'b0101001111;
    16'b0000100001001000: out_v[366] = 10'b0111000100;
    16'b1000100000001000: out_v[366] = 10'b1010110111;
    16'b0000100100000000: out_v[366] = 10'b0101111000;
    16'b1001100110001000: out_v[366] = 10'b1101010110;
    16'b0001100011001000: out_v[366] = 10'b0010110101;
    16'b0001100001101000: out_v[366] = 10'b0011101000;
    16'b0001100001001000: out_v[366] = 10'b1010001000;
    16'b0001100000101000: out_v[366] = 10'b1100011010;
    16'b0000100101100000: out_v[366] = 10'b1001011100;
    16'b0000100001100000: out_v[366] = 10'b1010010010;
    16'b0001100101100000: out_v[366] = 10'b0010010001;
    16'b1001100001001000: out_v[366] = 10'b1101001111;
    16'b0001100111001000: out_v[366] = 10'b0111101001;
    16'b0001100101101000: out_v[366] = 10'b1010000100;
    16'b0001100001100000: out_v[366] = 10'b0011010110;
    16'b0001100101000000: out_v[366] = 10'b0000111010;
    16'b0001100101100011: out_v[366] = 10'b1010011001;
    16'b1001100001101000: out_v[366] = 10'b0010100111;
    16'b0001100101101011: out_v[366] = 10'b1100000110;
    16'b0001100001100011: out_v[366] = 10'b0111000010;
    16'b0001100100001000: out_v[366] = 10'b0011011011;
    16'b0000000100100000: out_v[366] = 10'b0101000011;
    16'b0001100001000000: out_v[366] = 10'b0011101010;
    16'b0000100000100000: out_v[366] = 10'b0100111101;
    16'b0000100001100011: out_v[366] = 10'b0011010100;
    16'b1001100000001000: out_v[366] = 10'b1011111101;
    16'b0001000101101000: out_v[366] = 10'b0011011100;
    16'b0001100000001000: out_v[366] = 10'b1001100110;
    16'b1001100011001000: out_v[366] = 10'b0011111110;
    16'b0000100101100011: out_v[366] = 10'b1101100110;
    16'b0001100000100000: out_v[366] = 10'b0011011101;
    16'b0001000100101000: out_v[366] = 10'b1111100110;
    16'b0001100100101000: out_v[366] = 10'b0011101001;
    16'b1000000100000000: out_v[366] = 10'b1011101100;
    16'b0000000000100000: out_v[366] = 10'b1000011010;
    16'b1000100101001000: out_v[366] = 10'b0001111000;
    16'b1000000100101001: out_v[366] = 10'b1000111110;
    16'b1000000101001000: out_v[366] = 10'b0011001011;
    16'b1000000000001000: out_v[366] = 10'b0011011000;
    16'b1000000100001000: out_v[366] = 10'b0011011101;
    16'b0000000100100011: out_v[366] = 10'b0010101010;
    16'b0000000001000000: out_v[366] = 10'b1111011100;
    16'b0000000100100001: out_v[366] = 10'b0100111011;
    16'b0001000100000000: out_v[366] = 10'b0000111011;
    16'b0000000100101001: out_v[366] = 10'b0111110010;
    16'b1001000100001000: out_v[366] = 10'b1111010110;
    16'b1000100001001000: out_v[366] = 10'b0010011010;
    16'b0001000100100001: out_v[366] = 10'b1001110100;
    16'b0001000100101001: out_v[366] = 10'b0100010001;
    16'b0001000100101011: out_v[366] = 10'b0111001010;
    16'b1000000100101011: out_v[366] = 10'b0001011111;
    16'b1000000100101000: out_v[366] = 10'b0010011001;
    16'b0001000100100000: out_v[366] = 10'b0110011101;
    16'b0001000100100011: out_v[366] = 10'b0101001010;
    16'b1000000000000000: out_v[366] = 10'b0000101011;
    16'b1000000001001000: out_v[366] = 10'b0101011110;
    16'b0000000100101000: out_v[366] = 10'b0111110010;
    16'b0000100100100000: out_v[366] = 10'b0111100000;
    16'b0000100111000000: out_v[366] = 10'b1101001110;
    16'b0000100110001000: out_v[366] = 10'b0011011001;
    16'b0000100111001000: out_v[366] = 10'b1111001110;
    16'b0000100101001001: out_v[366] = 10'b1001110111;
    16'b0000100101000011: out_v[366] = 10'b0010110000;
    16'b0000100101000001: out_v[366] = 10'b1001010100;
    16'b0000110101000000: out_v[366] = 10'b0110011011;
    16'b0000100110000000: out_v[366] = 10'b1001110001;
    16'b0000100001000011: out_v[366] = 10'b0110110011;
    16'b0000100101001011: out_v[366] = 10'b0101101011;
    16'b0000100011001000: out_v[366] = 10'b0111100101;
    16'b0000100011000000: out_v[366] = 10'b0011011100;
    16'b0001000010001000: out_v[366] = 10'b0000110011;
    16'b0001000101000000: out_v[366] = 10'b1110100010;
    16'b1000100111001000: out_v[366] = 10'b1100101100;
    16'b0001000110001000: out_v[366] = 10'b0111011110;
    16'b1000000110001000: out_v[366] = 10'b1001001011;
    16'b0001000111001000: out_v[366] = 10'b1110100011;
    16'b0001100100000000: out_v[366] = 10'b1101011001;
    16'b0001000011001000: out_v[366] = 10'b1110111010;
    16'b0000000110001000: out_v[366] = 10'b0111000101;
    16'b1001000110001000: out_v[366] = 10'b0010010110;
    16'b0000000111001000: out_v[366] = 10'b1011101011;
    16'b0000000100101011: out_v[366] = 10'b0010100110;
    16'b0000000110101000: out_v[366] = 10'b1010011010;
    16'b0000110101100011: out_v[366] = 10'b0111011111;
    16'b0000100101100001: out_v[366] = 10'b1111000001;
    16'b0000100100100001: out_v[366] = 10'b1110110110;
    16'b0000110001100010: out_v[366] = 10'b0111101111;
    16'b0000110001100011: out_v[366] = 10'b0101101111;
    16'b0000000100000001: out_v[366] = 10'b1110000111;
    16'b0001110000100011: out_v[366] = 10'b1001011010;
    16'b0001110001100011: out_v[366] = 10'b1110100111;
    16'b0000100001100001: out_v[366] = 10'b1011001101;
    16'b0000010100100011: out_v[366] = 10'b1011010110;
    16'b0000100100100011: out_v[366] = 10'b1100000101;
    16'b0001110101100011: out_v[366] = 10'b1011011000;
    16'b0000100100000001: out_v[366] = 10'b1010101010;
    16'b0000110000100011: out_v[366] = 10'b1101100001;
    16'b0001100000100011: out_v[366] = 10'b1001110011;
    16'b0000100001000001: out_v[366] = 10'b0100010111;
    16'b0000100000100001: out_v[366] = 10'b0001111111;
    16'b0000100000100011: out_v[366] = 10'b1000010010;
    16'b0001110001000001: out_v[366] = 10'b1001000100;
    16'b1000100000000000: out_v[366] = 10'b0110011001;
    16'b1000100001000000: out_v[366] = 10'b1011101000;
    16'b1001100100001000: out_v[366] = 10'b0101110100;
    16'b0000000001001000: out_v[366] = 10'b0110100001;
    16'b1001100101001000: out_v[366] = 10'b0011100010;
    default: out_v[366] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000010000000: out_v[367] = 10'b1101001110;
    16'b0100000010000010: out_v[367] = 10'b1100001111;
    16'b0100000010000000: out_v[367] = 10'b0110011001;
    16'b0000000000000000: out_v[367] = 10'b1001100110;
    16'b0100000000000000: out_v[367] = 10'b1000100001;
    16'b0000010000000000: out_v[367] = 10'b1000011011;
    16'b0000010010000000: out_v[367] = 10'b0001100101;
    16'b0000000010000100: out_v[367] = 10'b0100011000;
    16'b0000000010000010: out_v[367] = 10'b1101001000;
    16'b0101000000000000: out_v[367] = 10'b1011110101;
    16'b0000000000000100: out_v[367] = 10'b1101110010;
    16'b0101000010000000: out_v[367] = 10'b1001001110;
    16'b0100000000000010: out_v[367] = 10'b0001100001;
    16'b0001000010000000: out_v[367] = 10'b0000100101;
    16'b0000010010000100: out_v[367] = 10'b1011110011;
    16'b0100010010000000: out_v[367] = 10'b0010111011;
    16'b0000010000000010: out_v[367] = 10'b1010011001;
    16'b0000010001000000: out_v[367] = 10'b1110010010;
    16'b0000010001000100: out_v[367] = 10'b1001100101;
    16'b0000010000000100: out_v[367] = 10'b1000011100;
    16'b0000010001001000: out_v[367] = 10'b0001000111;
    16'b0000000011000000: out_v[367] = 10'b0011000111;
    16'b0000010001001100: out_v[367] = 10'b0000011000;
    16'b0000000000100000: out_v[367] = 10'b1111000110;
    16'b0000010000100000: out_v[367] = 10'b1101111100;
    16'b0000000001000000: out_v[367] = 10'b1111011000;
    16'b0001010000000000: out_v[367] = 10'b0100001010;
    16'b0000000011001000: out_v[367] = 10'b1001010111;
    16'b0001000000000000: out_v[367] = 10'b0000100101;
    16'b0000000001001000: out_v[367] = 10'b1110100001;
    16'b0000001000000000: out_v[367] = 10'b0110100111;
    16'b0000000001000100: out_v[367] = 10'b0101001110;
    16'b0001010010000000: out_v[367] = 10'b0110001001;
    16'b0000000001001100: out_v[367] = 10'b0100101010;
    16'b0000010001001010: out_v[367] = 10'b1101110100;
    16'b0000000000000010: out_v[367] = 10'b0010111110;
    16'b0000010011000000: out_v[367] = 10'b0111001010;
    16'b0001010000000010: out_v[367] = 10'b0110100011;
    16'b0000010011001000: out_v[367] = 10'b1001111010;
    16'b0000010001000010: out_v[367] = 10'b1111110000;
    16'b0000010010000010: out_v[367] = 10'b1011101011;
    16'b0100010000000000: out_v[367] = 10'b1101000000;
    16'b0000000011000100: out_v[367] = 10'b0000110111;
    16'b0100000000000100: out_v[367] = 10'b0001100110;
    16'b0000000010100000: out_v[367] = 10'b0001100110;
    16'b0000010010100000: out_v[367] = 10'b0011001001;
    16'b0000000010000001: out_v[367] = 10'b1000010110;
    16'b0000010000001000: out_v[367] = 10'b0110100001;
    16'b0000010000000001: out_v[367] = 10'b1001100110;
    16'b0100010010000010: out_v[367] = 10'b1010001110;
    16'b0000010010000001: out_v[367] = 10'b0010010101;
    16'b0000000010001000: out_v[367] = 10'b0100011011;
    16'b0000010010001000: out_v[367] = 10'b1111011000;
    16'b0000000000001000: out_v[367] = 10'b0111001101;
    16'b0000010010000101: out_v[367] = 10'b0010111110;
    16'b0100010000000010: out_v[367] = 10'b1111111110;
    default: out_v[367] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000000001000: out_v[368] = 10'b1010001101;
    16'b0001000000001000: out_v[368] = 10'b1100000111;
    16'b0001100000001000: out_v[368] = 10'b1100100001;
    16'b0000000000000000: out_v[368] = 10'b0010110010;
    16'b0001100000000000: out_v[368] = 10'b1101110110;
    16'b0000100000000000: out_v[368] = 10'b1101110001;
    16'b0101000000000000: out_v[368] = 10'b0010111110;
    16'b0001000000000000: out_v[368] = 10'b1111110001;
    16'b0001000001001000: out_v[368] = 10'b0000110101;
    16'b0001100000000100: out_v[368] = 10'b0000100011;
    16'b0001000000000010: out_v[368] = 10'b0011001101;
    16'b0001000010000000: out_v[368] = 10'b1101100001;
    16'b0000100000001000: out_v[368] = 10'b0110001011;
    16'b0001100000001010: out_v[368] = 10'b1001000011;
    16'b0101100000001010: out_v[368] = 10'b0101010011;
    16'b0001000110000000: out_v[368] = 10'b1010110100;
    16'b0001000010001000: out_v[368] = 10'b0100011011;
    16'b0000100010000000: out_v[368] = 10'b1110010111;
    16'b0000100000000010: out_v[368] = 10'b0011100001;
    16'b0001000000001010: out_v[368] = 10'b0011001011;
    16'b0101100000000010: out_v[368] = 10'b1110011011;
    16'b0001100110000000: out_v[368] = 10'b1101111011;
    16'b0100000000001000: out_v[368] = 10'b0001101010;
    16'b0000000001001000: out_v[368] = 10'b1100001000;
    16'b0001100010000000: out_v[368] = 10'b0101111110;
    16'b0001000000000100: out_v[368] = 10'b1010111000;
    16'b0101000000001010: out_v[368] = 10'b1101010111;
    16'b0001100000000010: out_v[368] = 10'b1000100011;
    16'b0101000000001000: out_v[368] = 10'b0111110100;
    16'b0000000011001000: out_v[368] = 10'b0110001101;
    16'b0000000001000000: out_v[368] = 10'b1111000011;
    16'b0000000111001000: out_v[368] = 10'b0110000011;
    16'b0100000000000000: out_v[368] = 10'b1000001010;
    16'b0100000001000000: out_v[368] = 10'b1001000101;
    16'b0100000001001000: out_v[368] = 10'b1011101011;
    16'b0000000001001010: out_v[368] = 10'b1011001010;
    16'b0000000001000010: out_v[368] = 10'b1100011110;
    16'b0000100001001000: out_v[368] = 10'b0000110110;
    16'b0101000001001010: out_v[368] = 10'b1010000101;
    16'b0001000011000000: out_v[368] = 10'b0011001100;
    16'b0100000001001010: out_v[368] = 10'b0100001111;
    16'b0101000001001000: out_v[368] = 10'b0110100001;
    16'b0001100001001000: out_v[368] = 10'b1001101101;
    16'b0101100001001000: out_v[368] = 10'b0000011010;
    16'b0001000001001010: out_v[368] = 10'b0100011010;
    16'b0101000001000000: out_v[368] = 10'b1000110101;
    16'b0000000000001010: out_v[368] = 10'b1010111100;
    16'b0001000001000000: out_v[368] = 10'b1111000110;
    16'b0001000111001000: out_v[368] = 10'b1001001000;
    16'b0001000011001000: out_v[368] = 10'b1110001111;
    16'b0001100001000000: out_v[368] = 10'b0100011011;
    16'b0000100001000000: out_v[368] = 10'b1011100110;
    16'b0100000000001010: out_v[368] = 10'b0110111010;
    16'b0000000000000010: out_v[368] = 10'b1011010110;
    16'b0000000010001000: out_v[368] = 10'b0000011101;
    16'b0000000001000100: out_v[368] = 10'b1000111000;
    16'b0001100001001010: out_v[368] = 10'b1001011001;
    16'b0000000001001100: out_v[368] = 10'b1110010000;
    16'b0001100111001000: out_v[368] = 10'b0100011010;
    16'b0000100001001010: out_v[368] = 10'b1001111010;
    16'b0000000000000100: out_v[368] = 10'b0001110000;
    16'b0000000000001100: out_v[368] = 10'b1011100110;
    16'b0000000110000000: out_v[368] = 10'b1010100100;
    16'b0001000001001100: out_v[368] = 10'b1101011000;
    16'b0000000010000000: out_v[368] = 10'b0000110100;
    16'b0001000000001100: out_v[368] = 10'b1100010111;
    16'b0000000111000000: out_v[368] = 10'b0010111101;
    16'b0000000000000110: out_v[368] = 10'b1011110000;
    16'b0100000000000010: out_v[368] = 10'b1011110100;
    16'b0000000011000000: out_v[368] = 10'b1111001000;
    16'b0001000111000000: out_v[368] = 10'b1001001110;
    16'b0000001000001010: out_v[368] = 10'b0100011001;
    default: out_v[368] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010100000000100: out_v[369] = 10'b1100000110;
    16'b0100100010000111: out_v[369] = 10'b0100010000;
    16'b0101100010000111: out_v[369] = 10'b1100000111;
    16'b0001100000000100: out_v[369] = 10'b1100100110;
    16'b0100000010000011: out_v[369] = 10'b1100010111;
    16'b0100101110000111: out_v[369] = 10'b0000111111;
    16'b0101101110000111: out_v[369] = 10'b0000100001;
    16'b0000100000000100: out_v[369] = 10'b0011101110;
    16'b0100001110000011: out_v[369] = 10'b1111000111;
    16'b0100100010000110: out_v[369] = 10'b0001110101;
    16'b0111100010000111: out_v[369] = 10'b0110010101;
    16'b0110100010000111: out_v[369] = 10'b1110100010;
    16'b0011100000000100: out_v[369] = 10'b0011011000;
    16'b0000100000000101: out_v[369] = 10'b0110110001;
    16'b0100100010100111: out_v[369] = 10'b0001100101;
    16'b0100100000000100: out_v[369] = 10'b0011011011;
    16'b0100001110000111: out_v[369] = 10'b0111101010;
    16'b0000100000000000: out_v[369] = 10'b1100111011;
    16'b0101100000000100: out_v[369] = 10'b1101001011;
    16'b0100000010100011: out_v[369] = 10'b0011100001;
    16'b0100000010000010: out_v[369] = 10'b1001010101;
    16'b0111100000000101: out_v[369] = 10'b0110010010;
    16'b0100100000000101: out_v[369] = 10'b0011110111;
    16'b0101100000000101: out_v[369] = 10'b1101000011;
    16'b0100100010000011: out_v[369] = 10'b1110111111;
    16'b0010100000000101: out_v[369] = 10'b1101000111;
    16'b0101001110000111: out_v[369] = 10'b0010011110;
    16'b0000000010000011: out_v[369] = 10'b1001101100;
    16'b0111100010000110: out_v[369] = 10'b0101000011;
    16'b0100000010000111: out_v[369] = 10'b0010000011;
    16'b0000000000000000: out_v[369] = 10'b1101000011;
    16'b0000000000000001: out_v[369] = 10'b1000001111;
    16'b0000100010000111: out_v[369] = 10'b1011110011;
    16'b0101100010000110: out_v[369] = 10'b1011100111;
    16'b0111101110000111: out_v[369] = 10'b0101111111;
    16'b0100000010100111: out_v[369] = 10'b1011011100;
    16'b0001100010000111: out_v[369] = 10'b1110010100;
    16'b0110100000000101: out_v[369] = 10'b0010011011;
    16'b0010000000000100: out_v[369] = 10'b1001001111;
    16'b0000000000000100: out_v[369] = 10'b1100000011;
    16'b0000000000100000: out_v[369] = 10'b1001101010;
    16'b0000000000100001: out_v[369] = 10'b1011101100;
    16'b0010100000000000: out_v[369] = 10'b0111010111;
    16'b0010000000000000: out_v[369] = 10'b0110111110;
    16'b0001100000010100: out_v[369] = 10'b1011100000;
    16'b0000100000010100: out_v[369] = 10'b0101110100;
    16'b0001100001000100: out_v[369] = 10'b1010101010;
    16'b0001000001000100: out_v[369] = 10'b0000100100;
    16'b0001100000000101: out_v[369] = 10'b0101001101;
    16'b0000100010100111: out_v[369] = 10'b1011100101;
    16'b0001100000100101: out_v[369] = 10'b1001011100;
    16'b0001100000000000: out_v[369] = 10'b1111100110;
    16'b0101100011000110: out_v[369] = 10'b1011000101;
    16'b0000100001010100: out_v[369] = 10'b0010001111;
    16'b0000100010000110: out_v[369] = 10'b0000100000;
    16'b0001100010000110: out_v[369] = 10'b0100011010;
    16'b0001100001010100: out_v[369] = 10'b1010110111;
    16'b0100100010000010: out_v[369] = 10'b1010001100;
    16'b0001000000010100: out_v[369] = 10'b0011011101;
    16'b0001000000000000: out_v[369] = 10'b0011011010;
    16'b0000100000100100: out_v[369] = 10'b0111100100;
    16'b0001000001000000: out_v[369] = 10'b0100100110;
    16'b0000100000100101: out_v[369] = 10'b1001111110;
    16'b0100100011000110: out_v[369] = 10'b1111001100;
    16'b0001000000000100: out_v[369] = 10'b1110100001;
    16'b0001100000100100: out_v[369] = 10'b0010000101;
    16'b0011100000100100: out_v[369] = 10'b1110110011;
    16'b0011000000010100: out_v[369] = 10'b0001011110;
    16'b0011100000010100: out_v[369] = 10'b1100110110;
    16'b0011000000000100: out_v[369] = 10'b1110000101;
    16'b0011100000000101: out_v[369] = 10'b1001001011;
    16'b0011000000000000: out_v[369] = 10'b0010111101;
    16'b0000000000010100: out_v[369] = 10'b0111011001;
    16'b0100000000000001: out_v[369] = 10'b1001100100;
    16'b0100000000000000: out_v[369] = 10'b1010110100;
    16'b0101000010000010: out_v[369] = 10'b1110011010;
    16'b0100000000000101: out_v[369] = 10'b0001111011;
    16'b0101000010000011: out_v[369] = 10'b0011110010;
    16'b0011000000000001: out_v[369] = 10'b0000111110;
    16'b0000000000000101: out_v[369] = 10'b1000011011;
    16'b0111000000000001: out_v[369] = 10'b0101100111;
    16'b0101000000000000: out_v[369] = 10'b0010011111;
    16'b0001000000000001: out_v[369] = 10'b0111110010;
    16'b0111000000000000: out_v[369] = 10'b0110111111;
    16'b0110000000000000: out_v[369] = 10'b1101011101;
    16'b0101000000000001: out_v[369] = 10'b0101001010;
    16'b0110000000000001: out_v[369] = 10'b1101101111;
    16'b0110000010000011: out_v[369] = 10'b1011000100;
    16'b0100000010000110: out_v[369] = 10'b0000111010;
    16'b0111000010000011: out_v[369] = 10'b1010010111;
    16'b0010000000000001: out_v[369] = 10'b0110110001;
    16'b0110000010000010: out_v[369] = 10'b1101111010;
    16'b0000000010000110: out_v[369] = 10'b1010110010;
    16'b0000000010000010: out_v[369] = 10'b1000100110;
    16'b0010000000000101: out_v[369] = 10'b0111110100;
    16'b0011000000000101: out_v[369] = 10'b0100011100;
    16'b0100101110000110: out_v[369] = 10'b1111001110;
    16'b0101101110000110: out_v[369] = 10'b0111110110;
    16'b0101001100000000: out_v[369] = 10'b0110011001;
    16'b0101001110000010: out_v[369] = 10'b1101000011;
    16'b0001000000000101: out_v[369] = 10'b1110000011;
    16'b0101000000000100: out_v[369] = 10'b1000101011;
    16'b0100000000000100: out_v[369] = 10'b1010011111;
    16'b0101000010000110: out_v[369] = 10'b1010101000;
    16'b0110000000000101: out_v[369] = 10'b0011010110;
    16'b0110000010000111: out_v[369] = 10'b1101011010;
    16'b0101000010000111: out_v[369] = 10'b1000000111;
    16'b0110000000000100: out_v[369] = 10'b1001110110;
    default: out_v[369] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0101000001000000: out_v[370] = 10'b0110010101;
    16'b0101000000000000: out_v[370] = 10'b1001000011;
    16'b1101000000000000: out_v[370] = 10'b0101000100;
    16'b0000000000000000: out_v[370] = 10'b0001101011;
    16'b1001000000000000: out_v[370] = 10'b1000001001;
    16'b0001000000000000: out_v[370] = 10'b0001100011;
    16'b0101000100000000: out_v[370] = 10'b0110011110;
    16'b1101000001000000: out_v[370] = 10'b0011101110;
    16'b0100000000000000: out_v[370] = 10'b0110011011;
    16'b0101000000000010: out_v[370] = 10'b1010110010;
    16'b0101000001000010: out_v[370] = 10'b0111001001;
    16'b0001000001000000: out_v[370] = 10'b1000101010;
    16'b0100000001000000: out_v[370] = 10'b0011001000;
    16'b0001000000000010: out_v[370] = 10'b0100101110;
    16'b1100000000000000: out_v[370] = 10'b0100011101;
    16'b1101000000000010: out_v[370] = 10'b0100101011;
    16'b0001000000010000: out_v[370] = 10'b1101100001;
    16'b1101000001000010: out_v[370] = 10'b1111010011;
    16'b0000000100000000: out_v[370] = 10'b1011011100;
    16'b1000000100000000: out_v[370] = 10'b0101000110;
    16'b0000000101000000: out_v[370] = 10'b0011010111;
    16'b1000000101000000: out_v[370] = 10'b0011011010;
    16'b0001000100000000: out_v[370] = 10'b1101000010;
    16'b1001000100000000: out_v[370] = 10'b0000000111;
    16'b1000000000000000: out_v[370] = 10'b1000110101;
    16'b0101000100010000: out_v[370] = 10'b1110010011;
    16'b1101000100000000: out_v[370] = 10'b0111000100;
    16'b0000000100000010: out_v[370] = 10'b1011111101;
    16'b0100000100000010: out_v[370] = 10'b1111010000;
    16'b0101000100000010: out_v[370] = 10'b0011110111;
    16'b1001000100000010: out_v[370] = 10'b0011101110;
    16'b1100000100000000: out_v[370] = 10'b0100011111;
    16'b0100000100000000: out_v[370] = 10'b1000111100;
    16'b1101000100000010: out_v[370] = 10'b1010001100;
    16'b0001000100000010: out_v[370] = 10'b1101011110;
    16'b0101000101000000: out_v[370] = 10'b0001101100;
    16'b1101000101000000: out_v[370] = 10'b1110011011;
    16'b1001000101000000: out_v[370] = 10'b0111010100;
    16'b0000000001000000: out_v[370] = 10'b0010110011;
    16'b0100000101000010: out_v[370] = 10'b1111010001;
    16'b0000000101000010: out_v[370] = 10'b0101111000;
    16'b0001000101000000: out_v[370] = 10'b1000110001;
    16'b0001000101000010: out_v[370] = 10'b0011100111;
    16'b0101000101000010: out_v[370] = 10'b1100011010;
    16'b0001000001000010: out_v[370] = 10'b0000100111;
    16'b0100000101000000: out_v[370] = 10'b1001111000;
    16'b1001000001000000: out_v[370] = 10'b1001110111;
    16'b0000000001000010: out_v[370] = 10'b1000111110;
    16'b0111000100000000: out_v[370] = 10'b0111011100;
    16'b0110000100000000: out_v[370] = 10'b1011011111;
    16'b0100000100010000: out_v[370] = 10'b1110011010;
    16'b0011000000010000: out_v[370] = 10'b1011111111;
    16'b0011000100010000: out_v[370] = 10'b0000100010;
    16'b0011000100000000: out_v[370] = 10'b0011101010;
    16'b0001000100010000: out_v[370] = 10'b1001100000;
    16'b0011000000000000: out_v[370] = 10'b1010110110;
    16'b0100000001001010: out_v[370] = 10'b0101111010;
    16'b0100000100001000: out_v[370] = 10'b1010001111;
    16'b0100000001000010: out_v[370] = 10'b0111110111;
    16'b0100000000001010: out_v[370] = 10'b1101111110;
    16'b0100000000000010: out_v[370] = 10'b1011001000;
    16'b0100000100001010: out_v[370] = 10'b1101011111;
    16'b0100000000001000: out_v[370] = 10'b0001001100;
    16'b0000000100001010: out_v[370] = 10'b0101011001;
    16'b0000000000000010: out_v[370] = 10'b1011011101;
    16'b0000000100001000: out_v[370] = 10'b1001000111;
    default: out_v[370] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000010100000000: out_v[371] = 10'b1010100111;
    16'b0010010010000110: out_v[371] = 10'b1001000111;
    16'b0010010010000100: out_v[371] = 10'b1100110010;
    16'b1010010010000110: out_v[371] = 10'b0011011101;
    16'b0000010000000000: out_v[371] = 10'b0001011001;
    16'b1010000010000010: out_v[371] = 10'b1010111110;
    16'b0000010010000000: out_v[371] = 10'b0010000111;
    16'b0010000010000000: out_v[371] = 10'b1000100101;
    16'b1000010010000110: out_v[371] = 10'b0000011101;
    16'b0010000000000000: out_v[371] = 10'b0111000111;
    16'b0000010110000010: out_v[371] = 10'b1000101111;
    16'b0010010000000000: out_v[371] = 10'b1110001101;
    16'b0010000010000010: out_v[371] = 10'b0000111110;
    16'b0000010010000010: out_v[371] = 10'b1011110101;
    16'b0010010010000000: out_v[371] = 10'b1011010010;
    16'b0000010110000000: out_v[371] = 10'b0001001001;
    16'b0010000010000100: out_v[371] = 10'b1100010001;
    16'b0010010010000010: out_v[371] = 10'b1011000001;
    16'b1010000010000110: out_v[371] = 10'b1100000011;
    16'b1000010010000000: out_v[371] = 10'b0010110011;
    16'b0000000010000000: out_v[371] = 10'b1011100011;
    16'b0000010010000100: out_v[371] = 10'b0011001111;
    16'b0000010110000110: out_v[371] = 10'b1110110010;
    16'b0000010010000110: out_v[371] = 10'b0011010110;
    16'b1010010010000010: out_v[371] = 10'b1101011110;
    16'b0010000010000110: out_v[371] = 10'b0010101011;
    16'b1000010010000010: out_v[371] = 10'b1110000011;
    16'b0000010110000100: out_v[371] = 10'b1111010101;
    16'b0010000000000010: out_v[371] = 10'b1101011000;
    16'b0000000110000000: out_v[371] = 10'b0010010001;
    16'b0000010000000010: out_v[371] = 10'b0111100101;
    16'b0010010000000010: out_v[371] = 10'b0110011101;
    16'b1000010110000010: out_v[371] = 10'b1000011111;
    16'b1100000000000110: out_v[371] = 10'b0000001010;
    16'b0100000000000000: out_v[371] = 10'b1010010001;
    16'b0100010000000000: out_v[371] = 10'b0100011100;
    16'b0000000000000000: out_v[371] = 10'b0011001010;
    16'b1000000000000000: out_v[371] = 10'b0010111111;
    16'b0110010000000000: out_v[371] = 10'b0010010011;
    16'b1000000000000110: out_v[371] = 10'b1110110000;
    16'b1000000000000010: out_v[371] = 10'b0110011001;
    16'b0100000000000010: out_v[371] = 10'b1000011111;
    16'b0110000000000000: out_v[371] = 10'b1000001100;
    16'b1100000000000000: out_v[371] = 10'b0001110011;
    16'b0110010100000000: out_v[371] = 10'b1010100010;
    16'b1100000000000010: out_v[371] = 10'b1110100010;
    16'b0000000000000010: out_v[371] = 10'b0110011001;
    16'b0010010100000000: out_v[371] = 10'b0110001100;
    16'b0100000000000111: out_v[371] = 10'b1011100001;
    16'b0000000000000110: out_v[371] = 10'b0111110110;
    16'b0100000000000110: out_v[371] = 10'b0110000000;
    16'b0100010100000000: out_v[371] = 10'b0001001100;
    16'b0110000010000000: out_v[371] = 10'b0011010110;
    16'b1110000010000000: out_v[371] = 10'b0011000000;
    16'b1110000010000110: out_v[371] = 10'b1011100111;
    16'b0100000010000000: out_v[371] = 10'b1101100100;
    16'b1110000000000110: out_v[371] = 10'b1011001101;
    16'b1110000010000010: out_v[371] = 10'b0100110101;
    16'b0110000000000100: out_v[371] = 10'b0100111000;
    16'b0110000010000010: out_v[371] = 10'b1011001110;
    16'b0110000100000000: out_v[371] = 10'b0110011001;
    16'b0100010000000100: out_v[371] = 10'b0011100011;
    16'b0110000010000100: out_v[371] = 10'b0011110110;
    16'b1100010000000110: out_v[371] = 10'b0110000010;
    16'b0110010010000000: out_v[371] = 10'b0011011100;
    16'b0010000000000100: out_v[371] = 10'b1001111110;
    16'b1010000000000110: out_v[371] = 10'b1001110100;
    16'b0000010000000100: out_v[371] = 10'b1111011010;
    16'b0100010100000100: out_v[371] = 10'b1011011111;
    16'b0100010010000000: out_v[371] = 10'b1111100101;
    16'b0110000000000111: out_v[371] = 10'b1101100010;
    16'b1110010000000110: out_v[371] = 10'b0101011011;
    16'b0110010000000010: out_v[371] = 10'b0111110000;
    16'b0100000100000000: out_v[371] = 10'b0100000110;
    16'b0010010000000100: out_v[371] = 10'b1010100110;
    16'b0110010000000100: out_v[371] = 10'b1101110011;
    16'b0100010000000110: out_v[371] = 10'b0000011111;
    16'b0010010000000110: out_v[371] = 10'b1101100010;
    16'b1000010000000110: out_v[371] = 10'b1101011111;
    16'b0110010000000110: out_v[371] = 10'b0110110011;
    16'b0100010100000110: out_v[371] = 10'b1011111111;
    16'b0110000000000110: out_v[371] = 10'b0001011111;
    16'b0110010000000011: out_v[371] = 10'b0101001111;
    16'b1010010000000110: out_v[371] = 10'b1011110100;
    16'b0110010000000111: out_v[371] = 10'b1110001001;
    16'b0100010110000000: out_v[371] = 10'b1101101010;
    16'b0010000100000000: out_v[371] = 10'b0100011000;
    16'b0000000100000000: out_v[371] = 10'b1101000001;
    16'b0100010000000111: out_v[371] = 10'b1101011111;
    16'b0000010100000100: out_v[371] = 10'b0001110011;
    16'b0100000010000010: out_v[371] = 10'b0001011110;
    16'b0110000110000000: out_v[371] = 10'b0010111001;
    16'b0110000000100000: out_v[371] = 10'b0000110011;
    16'b0110000000000010: out_v[371] = 10'b0101100101;
    16'b0110010010000010: out_v[371] = 10'b0010110000;
    16'b1110010010000010: out_v[371] = 10'b1001010110;
    16'b0100000110000000: out_v[371] = 10'b1000011010;
    16'b0110010110000000: out_v[371] = 10'b0100110111;
    16'b0110000100000010: out_v[371] = 10'b0101110000;
    16'b0100000000100000: out_v[371] = 10'b1000001101;
    16'b1110010000000000: out_v[371] = 10'b1011110000;
    16'b0110000110000010: out_v[371] = 10'b0010000101;
    16'b0110010100000010: out_v[371] = 10'b0100011011;
    16'b0100000010100000: out_v[371] = 10'b0101111010;
    16'b0110000010100000: out_v[371] = 10'b0010011011;
    16'b0110010010100000: out_v[371] = 10'b0010010010;
    16'b0110010110000010: out_v[371] = 10'b0010011001;
    16'b0100010100000010: out_v[371] = 10'b1000100110;
    16'b0010010000100110: out_v[371] = 10'b0011011110;
    16'b0100000100000010: out_v[371] = 10'b0001110111;
    16'b0110010000100110: out_v[371] = 10'b1111001010;
    16'b1000010000000000: out_v[371] = 10'b1010111010;
    16'b1100010100000010: out_v[371] = 10'b1000110111;
    16'b1110010000000010: out_v[371] = 10'b1010100000;
    16'b0110010000100010: out_v[371] = 10'b0111001110;
    16'b0010010000100010: out_v[371] = 10'b1011111111;
    16'b0010010100000010: out_v[371] = 10'b1110111100;
    16'b1100010100000000: out_v[371] = 10'b0010100111;
    16'b0100010000000010: out_v[371] = 10'b0110000000;
    16'b0000010100000010: out_v[371] = 10'b0011100110;
    16'b0010010100100010: out_v[371] = 10'b1010111011;
    16'b1100010000000010: out_v[371] = 10'b1110100101;
    16'b1100010000000000: out_v[371] = 10'b0110110110;
    16'b1110010010000000: out_v[371] = 10'b1110100010;
    16'b1110000000000000: out_v[371] = 10'b0011110010;
    16'b1010000000000000: out_v[371] = 10'b1001100000;
    16'b1010010000000000: out_v[371] = 10'b1101011001;
    16'b1010000010000000: out_v[371] = 10'b1001100110;
    16'b1100010010000010: out_v[371] = 10'b1001111001;
    16'b1010010000000010: out_v[371] = 10'b1001001001;
    16'b1100000010000000: out_v[371] = 10'b0111010111;
    16'b1110000000000010: out_v[371] = 10'b1110100011;
    16'b1100010010000000: out_v[371] = 10'b1011011011;
    16'b0111000100000000: out_v[371] = 10'b1101101111;
    16'b0011010000000000: out_v[371] = 10'b1110101011;
    16'b0001000100000000: out_v[371] = 10'b1010100110;
    16'b0111010100000000: out_v[371] = 10'b1100000101;
    16'b0111010000000000: out_v[371] = 10'b1010100111;
    16'b0110000000000001: out_v[371] = 10'b0101011010;
    16'b0100000000000101: out_v[371] = 10'b0011110000;
    16'b0100000000000001: out_v[371] = 10'b1010000111;
    16'b0011010100000000: out_v[371] = 10'b1100111010;
    16'b0011000100000000: out_v[371] = 10'b0101101110;
    16'b0110010010000110: out_v[371] = 10'b1110111110;
    16'b0110010000100000: out_v[371] = 10'b0111001111;
    16'b0010000110000000: out_v[371] = 10'b1110001110;
    16'b0101000100000000: out_v[371] = 10'b1101100111;
    default: out_v[371] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000100001001101: out_v[372] = 10'b1000011000;
    16'b0100100001001001: out_v[372] = 10'b1000000111;
    16'b0100100000001000: out_v[372] = 10'b1010101111;
    16'b0100000000010000: out_v[372] = 10'b0111100101;
    16'b0100100001001000: out_v[372] = 10'b1011001010;
    16'b0100000001000000: out_v[372] = 10'b0111100110;
    16'b0100000000000000: out_v[372] = 10'b0011010010;
    16'b0000100000001100: out_v[372] = 10'b0100001111;
    16'b0100100001001101: out_v[372] = 10'b1101101000;
    16'b0000100000001101: out_v[372] = 10'b0111011010;
    16'b0000000000001100: out_v[372] = 10'b1000011010;
    16'b0000100001001000: out_v[372] = 10'b1101011111;
    16'b0000100001001001: out_v[372] = 10'b0011111011;
    16'b0100100001001100: out_v[372] = 10'b0110100000;
    16'b0100100000001001: out_v[372] = 10'b1111000111;
    16'b0100000000001000: out_v[372] = 10'b0011111011;
    16'b0100100000001100: out_v[372] = 10'b0010110110;
    16'b0000100000001001: out_v[372] = 10'b1011000110;
    16'b0000000000000100: out_v[372] = 10'b1011101000;
    16'b0100000001000001: out_v[372] = 10'b0001000011;
    16'b0000100001001100: out_v[372] = 10'b1010101001;
    16'b0100100000001101: out_v[372] = 10'b1001001100;
    16'b0000100000011100: out_v[372] = 10'b0110100111;
    16'b0000000000000101: out_v[372] = 10'b1000111011;
    16'b0000100000001000: out_v[372] = 10'b0100000100;
    16'b0100000001001001: out_v[372] = 10'b1001110110;
    16'b0000000000001101: out_v[372] = 10'b0101010010;
    16'b0100100000011100: out_v[372] = 10'b1100101000;
    16'b0100000000001101: out_v[372] = 10'b0111010101;
    16'b0100100000011000: out_v[372] = 10'b1011111100;
    16'b0100000000000100: out_v[372] = 10'b0100011100;
    16'b0100000000001100: out_v[372] = 10'b0110100111;
    16'b0000000000000000: out_v[372] = 10'b1011101001;
    16'b0100100000000000: out_v[372] = 10'b0100011111;
    16'b0000100000000000: out_v[372] = 10'b0010000010;
    16'b0000000001000000: out_v[372] = 10'b0110011110;
    16'b0000000001010001: out_v[372] = 10'b0100100100;
    16'b0100000001001000: out_v[372] = 10'b1011100101;
    16'b0100100011001001: out_v[372] = 10'b1001011110;
    16'b0100100001011001: out_v[372] = 10'b0010010100;
    16'b0100000001010000: out_v[372] = 10'b1001110110;
    16'b0100100000011001: out_v[372] = 10'b1100100111;
    16'b0000100001011001: out_v[372] = 10'b0000111110;
    16'b0100100001011000: out_v[372] = 10'b0101010101;
    16'b0000000000000001: out_v[372] = 10'b0010101100;
    16'b0000000001000001: out_v[372] = 10'b1100010110;
    16'b0100000001010001: out_v[372] = 10'b1011111000;
    16'b0100000001011000: out_v[372] = 10'b1111011000;
    16'b0000000001010000: out_v[372] = 10'b1101000110;
    16'b0100000000011000: out_v[372] = 10'b1110011010;
    16'b0000000001001000: out_v[372] = 10'b1111010110;
    16'b0000000001000100: out_v[372] = 10'b1010011000;
    16'b0000000001001101: out_v[372] = 10'b0011010110;
    16'b0000000001001100: out_v[372] = 10'b0010101011;
    16'b0100100011001000: out_v[372] = 10'b0110010100;
    16'b0100000001000100: out_v[372] = 10'b0110110011;
    16'b0000000001000101: out_v[372] = 10'b1000110100;
    16'b0100000001001100: out_v[372] = 10'b0011011001;
    16'b0000000000001000: out_v[372] = 10'b0110110011;
    16'b0100100000000001: out_v[372] = 10'b0100111000;
    16'b0100000000000001: out_v[372] = 10'b0101011010;
    16'b0100000000000101: out_v[372] = 10'b1110001010;
    16'b0000100001000001: out_v[372] = 10'b0010110010;
    16'b0100000001000101: out_v[372] = 10'b0110110001;
    16'b0000000001001001: out_v[372] = 10'b0011010011;
    16'b0000100001000101: out_v[372] = 10'b0001011001;
    16'b0100100001000001: out_v[372] = 10'b1101010011;
    16'b0000100000000101: out_v[372] = 10'b0110110111;
    16'b0100000000010001: out_v[372] = 10'b1011000111;
    16'b0100000000001001: out_v[372] = 10'b0011110011;
    16'b0100000000100000: out_v[372] = 10'b1010000111;
    16'b0100000001100000: out_v[372] = 10'b0111011011;
    16'b0001000001000001: out_v[372] = 10'b1001101111;
    default: out_v[372] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010000000000000: out_v[373] = 10'b0010010110;
    16'b0011000000000000: out_v[373] = 10'b1100000001;
    16'b0001000000000000: out_v[373] = 10'b0001110100;
    16'b0000000000000000: out_v[373] = 10'b0100011000;
    16'b0110000000000000: out_v[373] = 10'b0000001111;
    16'b0100000000000000: out_v[373] = 10'b0101110100;
    16'b0111000000000000: out_v[373] = 10'b0001001111;
    16'b0101000000000000: out_v[373] = 10'b0101011011;
    16'b0011000000000100: out_v[373] = 10'b0100001001;
    16'b0000000000000010: out_v[373] = 10'b0000011110;
    16'b0000000010000000: out_v[373] = 10'b0101100000;
    16'b0010000000000010: out_v[373] = 10'b1110011011;
    16'b0010000000001000: out_v[373] = 10'b0010001000;
    16'b0010010000000000: out_v[373] = 10'b1000100101;
    16'b0000000000000100: out_v[373] = 10'b0000100001;
    16'b0000010000000000: out_v[373] = 10'b1100000000;
    16'b0010000000000100: out_v[373] = 10'b0100110000;
    16'b0000000000100000: out_v[373] = 10'b0000101000;
    16'b0010000000100000: out_v[373] = 10'b0101100100;
    16'b0010000000100100: out_v[373] = 10'b0010111100;
    16'b0000000100000000: out_v[373] = 10'b1001110001;
    16'b0010000100000000: out_v[373] = 10'b1101001011;
    16'b0001000010000000: out_v[373] = 10'b1111100111;
    16'b0100000010000000: out_v[373] = 10'b0011001111;
    16'b0010000000010000: out_v[373] = 10'b1000001000;
    16'b0000000000010000: out_v[373] = 10'b1011000101;
    16'b0011000000100000: out_v[373] = 10'b0111011101;
    16'b0001000000100000: out_v[373] = 10'b0010011010;
    default: out_v[373] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1000001010000000: out_v[374] = 10'b0100100001;
    16'b1000001010100000: out_v[374] = 10'b0111010101;
    16'b0000001000100000: out_v[374] = 10'b0010010110;
    16'b0000000010000000: out_v[374] = 10'b1101111000;
    16'b0000001010000000: out_v[374] = 10'b1100001001;
    16'b0000000000100000: out_v[374] = 10'b0101010001;
    16'b0010001000100000: out_v[374] = 10'b1010000101;
    16'b0000001010100000: out_v[374] = 10'b1001100100;
    16'b1010001010000000: out_v[374] = 10'b1101010010;
    16'b0000001000000000: out_v[374] = 10'b1000000110;
    16'b0000000000000000: out_v[374] = 10'b1000010110;
    16'b0000000010100000: out_v[374] = 10'b0111010011;
    16'b1000000010000000: out_v[374] = 10'b0010011111;
    16'b0010001010100000: out_v[374] = 10'b0000010011;
    16'b1010001010100000: out_v[374] = 10'b0100111100;
    16'b0010001010000000: out_v[374] = 10'b0110001010;
    16'b1010001000000000: out_v[374] = 10'b0110001010;
    16'b0010001000000000: out_v[374] = 10'b0010001100;
    16'b1000001000000000: out_v[374] = 10'b0101101001;
    16'b1000000000000000: out_v[374] = 10'b1001001111;
    16'b0010000000000000: out_v[374] = 10'b1001001110;
    16'b1010000010000000: out_v[374] = 10'b0111010000;
    16'b1010000000000000: out_v[374] = 10'b1100000000;
    16'b1000000010100000: out_v[374] = 10'b0000110100;
    16'b1010000010100000: out_v[374] = 10'b1100101010;
    16'b0010000000100000: out_v[374] = 10'b1001110001;
    16'b1010001000100000: out_v[374] = 10'b0111010111;
    16'b0000001100000000: out_v[374] = 10'b0011011110;
    16'b1010001110000000: out_v[374] = 10'b1101011010;
    16'b1010001010100001: out_v[374] = 10'b1011111001;
    16'b1010000110000000: out_v[374] = 10'b0110010110;
    16'b1010001011100000: out_v[374] = 10'b0001011001;
    16'b1010001110100000: out_v[374] = 10'b1110100100;
    16'b0010000010000000: out_v[374] = 10'b0111010011;
    16'b0010000010100000: out_v[374] = 10'b1001110010;
    16'b1010000000100000: out_v[374] = 10'b0011001000;
    16'b0000001000010000: out_v[374] = 10'b0011110110;
    16'b0010001001000000: out_v[374] = 10'b1010110111;
    16'b0000001001000000: out_v[374] = 10'b1111110110;
    16'b0010011000000000: out_v[374] = 10'b1101100101;
    default: out_v[374] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010000101000000: out_v[375] = 10'b1100010010;
    16'b1110000001000000: out_v[375] = 10'b0001111011;
    16'b0110000101100000: out_v[375] = 10'b1000100011;
    16'b1110000101100000: out_v[375] = 10'b1011110101;
    16'b0110000101000000: out_v[375] = 10'b0010000011;
    16'b0010000101100000: out_v[375] = 10'b1100010001;
    16'b0100000101100000: out_v[375] = 10'b0011111101;
    16'b0000000100100000: out_v[375] = 10'b0000111100;
    16'b0110100101100000: out_v[375] = 10'b1011111000;
    16'b0010000100100000: out_v[375] = 10'b1110010111;
    16'b0000000100000000: out_v[375] = 10'b0010110001;
    16'b0010000100000000: out_v[375] = 10'b1010100001;
    16'b1110000101000000: out_v[375] = 10'b0110100100;
    16'b0110000100000000: out_v[375] = 10'b0011110111;
    16'b0000000000100000: out_v[375] = 10'b0101110011;
    16'b1010000100100000: out_v[375] = 10'b0001010111;
    16'b0010000001000000: out_v[375] = 10'b0101110000;
    16'b1110000001100000: out_v[375] = 10'b0010111111;
    16'b1010000101100000: out_v[375] = 10'b1110110011;
    16'b0000000101000000: out_v[375] = 10'b1100110011;
    16'b0000000000000000: out_v[375] = 10'b0010010101;
    16'b0110000100100000: out_v[375] = 10'b0100001011;
    16'b0110000001000000: out_v[375] = 10'b0001011111;
    16'b1010000101000000: out_v[375] = 10'b1110110011;
    16'b0100000001100000: out_v[375] = 10'b1101000100;
    16'b0100000001000000: out_v[375] = 10'b0010010110;
    16'b1110100101100000: out_v[375] = 10'b0010001001;
    16'b1010100100100000: out_v[375] = 10'b1101111001;
    16'b0100000000100000: out_v[375] = 10'b0011110010;
    16'b1010000100000000: out_v[375] = 10'b1010101001;
    16'b1000000000000000: out_v[375] = 10'b0010011011;
    16'b0100000000000000: out_v[375] = 10'b1011000011;
    16'b0110000000000000: out_v[375] = 10'b1000011010;
    16'b1000010000000000: out_v[375] = 10'b0110111010;
    16'b0000000001000000: out_v[375] = 10'b0001001100;
    16'b0100000001000010: out_v[375] = 10'b0101000100;
    16'b1100000000000000: out_v[375] = 10'b0010111111;
    16'b0100000000000010: out_v[375] = 10'b1110100011;
    16'b0100100001000000: out_v[375] = 10'b0011001011;
    16'b0000100000000000: out_v[375] = 10'b1001111100;
    16'b0000000001000010: out_v[375] = 10'b1010111100;
    16'b1100000001000000: out_v[375] = 10'b0000001000;
    16'b0000100001000000: out_v[375] = 10'b0000110110;
    16'b0001000001000000: out_v[375] = 10'b1001010101;
    16'b1000000001000000: out_v[375] = 10'b0010001001;
    16'b0101000001000000: out_v[375] = 10'b0011010111;
    16'b0011000101000000: out_v[375] = 10'b0110111100;
    16'b0100000101000000: out_v[375] = 10'b1110100011;
    16'b1110000100000000: out_v[375] = 10'b0100001110;
    16'b0001000000000000: out_v[375] = 10'b1110101011;
    16'b0010100101000000: out_v[375] = 10'b0111100101;
    16'b1010000000000000: out_v[375] = 10'b1100011010;
    16'b1000100001000000: out_v[375] = 10'b1100110010;
    16'b0010000000000000: out_v[375] = 10'b1101011001;
    16'b1100100001000000: out_v[375] = 10'b0001000011;
    16'b1010000001000000: out_v[375] = 10'b0001101111;
    16'b1000100000000000: out_v[375] = 10'b0111001011;
    16'b0010000111000000: out_v[375] = 10'b1010100000;
    16'b0100000100000000: out_v[375] = 10'b1101111000;
    16'b0010010100000000: out_v[375] = 10'b1101000000;
    16'b0010010000000000: out_v[375] = 10'b1110101100;
    16'b0000000111000000: out_v[375] = 10'b0010101101;
    16'b0000000011000000: out_v[375] = 10'b1101001000;
    16'b0110010100000000: out_v[375] = 10'b0110000110;
    16'b0110010101000000: out_v[375] = 10'b1011110110;
    16'b0010010101000000: out_v[375] = 10'b1000101000;
    16'b1110010101000000: out_v[375] = 10'b0110110000;
    16'b0110010001000000: out_v[375] = 10'b0110101111;
    16'b1110010100000000: out_v[375] = 10'b0011100011;
    16'b1010010101000000: out_v[375] = 10'b1101010011;
    16'b0100010001000000: out_v[375] = 10'b0000000011;
    16'b0110000101001000: out_v[375] = 10'b1011000010;
    16'b0100000001100010: out_v[375] = 10'b1111101111;
    16'b0100000101001000: out_v[375] = 10'b1101101010;
    16'b0010000101000001: out_v[375] = 10'b1111101111;
    16'b0110000111000000: out_v[375] = 10'b0111110111;
    16'b0010000111000001: out_v[375] = 10'b0110010011;
    16'b1110000100100000: out_v[375] = 10'b0101101011;
    16'b1010010100000000: out_v[375] = 10'b1011101110;
    16'b1110000000000000: out_v[375] = 10'b1101110011;
    default: out_v[375] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001000000000001: out_v[376] = 10'b0011010011;
    16'b0000000000000011: out_v[376] = 10'b0001001010;
    16'b0001000001000000: out_v[376] = 10'b0100100111;
    16'b0001000000010111: out_v[376] = 10'b1101101110;
    16'b0000000000000001: out_v[376] = 10'b0100011111;
    16'b0001000000000000: out_v[376] = 10'b1010111100;
    16'b0000000000010000: out_v[376] = 10'b1010101001;
    16'b0000000000000000: out_v[376] = 10'b1010100100;
    16'b0001000001000011: out_v[376] = 10'b0110011101;
    16'b0000000001000000: out_v[376] = 10'b0100100101;
    16'b0000000000010011: out_v[376] = 10'b1100001111;
    16'b0001000000000101: out_v[376] = 10'b1100100010;
    16'b0001000000000100: out_v[376] = 10'b1001011011;
    16'b0001000000010001: out_v[376] = 10'b1011010110;
    16'b0000000000000101: out_v[376] = 10'b1100001101;
    16'b0001000000010101: out_v[376] = 10'b1001001111;
    16'b0000000000000010: out_v[376] = 10'b0000011111;
    16'b0001000001000111: out_v[376] = 10'b0100110011;
    16'b0001000001000101: out_v[376] = 10'b1111010010;
    16'b0001000010000101: out_v[376] = 10'b0000101011;
    16'b0001000000010011: out_v[376] = 10'b1000001100;
    16'b0001000000000011: out_v[376] = 10'b0101010000;
    16'b0000000100000010: out_v[376] = 10'b0110001011;
    16'b0000000001000010: out_v[376] = 10'b0110010011;
    16'b0001000001000100: out_v[376] = 10'b1111010000;
    16'b0000000100010010: out_v[376] = 10'b0110000101;
    16'b0000000100000011: out_v[376] = 10'b1101100100;
    16'b0001000100010011: out_v[376] = 10'b1100000111;
    16'b0001000001000001: out_v[376] = 10'b1110001111;
    16'b0001000000010000: out_v[376] = 10'b1011000101;
    16'b0000000000010010: out_v[376] = 10'b1111110000;
    16'b0001000000000111: out_v[376] = 10'b1011101110;
    16'b0000000001000011: out_v[376] = 10'b1001011011;
    16'b0001000000000010: out_v[376] = 10'b1001110010;
    16'b0000000100010011: out_v[376] = 10'b1011111011;
    16'b0000000000010001: out_v[376] = 10'b0101010111;
    16'b0000000000000100: out_v[376] = 10'b0110110100;
    16'b0000000010000101: out_v[376] = 10'b0010101101;
    16'b0000000010000001: out_v[376] = 10'b0101001110;
    16'b1001000010000101: out_v[376] = 10'b0111110010;
    16'b0001000010000001: out_v[376] = 10'b0100001101;
    16'b0001000010000111: out_v[376] = 10'b0100110101;
    16'b0001000100000011: out_v[376] = 10'b1111010101;
    16'b0001000100000111: out_v[376] = 10'b0001000011;
    16'b0001000010000100: out_v[376] = 10'b0000100110;
    16'b0000000010000100: out_v[376] = 10'b1001100101;
    16'b0000000000000111: out_v[376] = 10'b1001101110;
    16'b0000010000000000: out_v[376] = 10'b1010001000;
    16'b0001000110000101: out_v[376] = 10'b1100011110;
    16'b0000000100000101: out_v[376] = 10'b0101001011;
    16'b0001010000000100: out_v[376] = 10'b1001001010;
    16'b0000000100000001: out_v[376] = 10'b0111110011;
    16'b0000010000000100: out_v[376] = 10'b0100011011;
    16'b0001000100000101: out_v[376] = 10'b0011001001;
    16'b0001000110000111: out_v[376] = 10'b0011100111;
    16'b0000000100000111: out_v[376] = 10'b1000100100;
    16'b0001000010000000: out_v[376] = 10'b0001111100;
    16'b0000000010000000: out_v[376] = 10'b1111010000;
    16'b0000000000000110: out_v[376] = 10'b1000010001;
    16'b0001000000010010: out_v[376] = 10'b0000010110;
    16'b0000000100000000: out_v[376] = 10'b0111011010;
    16'b0001000000000110: out_v[376] = 10'b1010110010;
    16'b0000000001000001: out_v[376] = 10'b0011100110;
    16'b0001000000001000: out_v[376] = 10'b1010101000;
    16'b0000000000001000: out_v[376] = 10'b1010000000;
    16'b0000010001000000: out_v[376] = 10'b1011011110;
    default: out_v[376] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0100010000100000: out_v[377] = 10'b0011101010;
    16'b0100111000000000: out_v[377] = 10'b0010010111;
    16'b0100110000000000: out_v[377] = 10'b0101101011;
    16'b0000110000100000: out_v[377] = 10'b1010010000;
    16'b0110100000110000: out_v[377] = 10'b0000110111;
    16'b0100111000100001: out_v[377] = 10'b1000011011;
    16'b0100001000000001: out_v[377] = 10'b1110101111;
    16'b0100100000000000: out_v[377] = 10'b0101011011;
    16'b0100001000010000: out_v[377] = 10'b1011001011;
    16'b0010110000100000: out_v[377] = 10'b0001111000;
    16'b0100111000000001: out_v[377] = 10'b0000101011;
    16'b0000111000000001: out_v[377] = 10'b0011111001;
    16'b0000011000000000: out_v[377] = 10'b1100011111;
    16'b0100011000000100: out_v[377] = 10'b0111111101;
    16'b0100000000010000: out_v[377] = 10'b1011000001;
    16'b0100011000000000: out_v[377] = 10'b1001100110;
    16'b0100011000000001: out_v[377] = 10'b1010110010;
    16'b0000111000000000: out_v[377] = 10'b0111001001;
    16'b0100101000010001: out_v[377] = 10'b1111011011;
    16'b0110110000110000: out_v[377] = 10'b1010111001;
    16'b0100100000010000: out_v[377] = 10'b1000001010;
    16'b0100101000010000: out_v[377] = 10'b0100110111;
    16'b0000100000010000: out_v[377] = 10'b0011110101;
    16'b0100111000010001: out_v[377] = 10'b0111011110;
    16'b0100001000010101: out_v[377] = 10'b1010101110;
    16'b0100001000010100: out_v[377] = 10'b1111010111;
    16'b0000111000100000: out_v[377] = 10'b1010000010;
    16'b0100101000000000: out_v[377] = 10'b0011110110;
    16'b0100101000000001: out_v[377] = 10'b1111000110;
    16'b0100100000110000: out_v[377] = 10'b0101001101;
    16'b0100110000110000: out_v[377] = 10'b1011010000;
    16'b0110111000100001: out_v[377] = 10'b0101010011;
    16'b0100001000000000: out_v[377] = 10'b0011001111;
    16'b0100100000010001: out_v[377] = 10'b1011111111;
    16'b0010111010000001: out_v[377] = 10'b1010010011;
    16'b0100110000000001: out_v[377] = 10'b0101101111;
    16'b0010111000000001: out_v[377] = 10'b1011000101;
    16'b0100110000100000: out_v[377] = 10'b1001000110;
    16'b0000111000100001: out_v[377] = 10'b0001011011;
    16'b0110111000000001: out_v[377] = 10'b1101011011;
    16'b0000010000100000: out_v[377] = 10'b1010000001;
    16'b0000000000010000: out_v[377] = 10'b1111000011;
    16'b0000110010100000: out_v[377] = 10'b1100011111;
    16'b0100000000010100: out_v[377] = 10'b0011001111;
    16'b0100010000000000: out_v[377] = 10'b0010111110;
    16'b0110110000100000: out_v[377] = 10'b1001110000;
    16'b0100001000010001: out_v[377] = 10'b0111001010;
    16'b0100111000100000: out_v[377] = 10'b0110110010;
    16'b0100000000010001: out_v[377] = 10'b1100011101;
    16'b0100000000000000: out_v[377] = 10'b1100100110;
    16'b0000110000000000: out_v[377] = 10'b1011001000;
    16'b0000010000000000: out_v[377] = 10'b1100101100;
    16'b0010100010100000: out_v[377] = 10'b1011110000;
    16'b0010100010100100: out_v[377] = 10'b1001110111;
    16'b0010000010000000: out_v[377] = 10'b0110010101;
    16'b0000100010000000: out_v[377] = 10'b0011001100;
    16'b0000000010000000: out_v[377] = 10'b1010100111;
    16'b0010100010000000: out_v[377] = 10'b0000111010;
    16'b0010000000000000: out_v[377] = 10'b1001000011;
    16'b0010101010100000: out_v[377] = 10'b1000001011;
    16'b0010100010000100: out_v[377] = 10'b0110000110;
    16'b0010001010100000: out_v[377] = 10'b0001010110;
    16'b0010101010000000: out_v[377] = 10'b0111001100;
    16'b0010001010000000: out_v[377] = 10'b0100010010;
    16'b0000000000000000: out_v[377] = 10'b0000100010;
    16'b0010100000000000: out_v[377] = 10'b1100010110;
    16'b0010100010010000: out_v[377] = 10'b1011010101;
    16'b0010100110010000: out_v[377] = 10'b1000011100;
    16'b0000110010000000: out_v[377] = 10'b1011100010;
    16'b0010100000010000: out_v[377] = 10'b0110010011;
    16'b0010100010110000: out_v[377] = 10'b0101011010;
    16'b0010100000110000: out_v[377] = 10'b0100101000;
    16'b0000110010110000: out_v[377] = 10'b0110010100;
    16'b0000111000010001: out_v[377] = 10'b1011110100;
    16'b0000111000110001: out_v[377] = 10'b1101010010;
    16'b0000111010010001: out_v[377] = 10'b0110010110;
    16'b0010110000000000: out_v[377] = 10'b0000010111;
    16'b0000110000110000: out_v[377] = 10'b1101110110;
    16'b0010110010000000: out_v[377] = 10'b1110100100;
    16'b0010110010110000: out_v[377] = 10'b0100101010;
    16'b0000110010100001: out_v[377] = 10'b0101110110;
    16'b0010100110110000: out_v[377] = 10'b0011111010;
    16'b0000101000110001: out_v[377] = 10'b0110100111;
    16'b0010010010000000: out_v[377] = 10'b0100001000;
    16'b0000110000100001: out_v[377] = 10'b0101100001;
    16'b0010110010100000: out_v[377] = 10'b1011000100;
    16'b0000100000110000: out_v[377] = 10'b0001101111;
    16'b0010101010110000: out_v[377] = 10'b1011110101;
    16'b0000111010100001: out_v[377] = 10'b1101101110;
    16'b0010100000100000: out_v[377] = 10'b1101101101;
    16'b0010110000110000: out_v[377] = 10'b1011101000;
    16'b0110110010000000: out_v[377] = 10'b0111100110;
    16'b0000111010110001: out_v[377] = 10'b1010111001;
    16'b0010110010010000: out_v[377] = 10'b1011001010;
    16'b0000100000100000: out_v[377] = 10'b0011100101;
    16'b0110110010100000: out_v[377] = 10'b1111100110;
    16'b0000111010000001: out_v[377] = 10'b1010010110;
    16'b0010000010010000: out_v[377] = 10'b1001001100;
    16'b0110100010010000: out_v[377] = 10'b0001110111;
    16'b0000101000100001: out_v[377] = 10'b1010110101;
    16'b0110100010110000: out_v[377] = 10'b1001001001;
    16'b0010010010100100: out_v[377] = 10'b1111110010;
    16'b0010111000100001: out_v[377] = 10'b1010111100;
    16'b0010110010100001: out_v[377] = 10'b1101101010;
    16'b0010010010100000: out_v[377] = 10'b1011100011;
    16'b0010010010000100: out_v[377] = 10'b0100100111;
    16'b0010010010010100: out_v[377] = 10'b1010100110;
    16'b0010010000100100: out_v[377] = 10'b0001001010;
    16'b0010010010100001: out_v[377] = 10'b1010101101;
    16'b0010000010000100: out_v[377] = 10'b0101001000;
    16'b0000000010010000: out_v[377] = 10'b1011001111;
    16'b0010000010010100: out_v[377] = 10'b1001110110;
    16'b0010000010100000: out_v[377] = 10'b0010111001;
    16'b0010111010100001: out_v[377] = 10'b1001001010;
    16'b0010000010110100: out_v[377] = 10'b0110011011;
    16'b0000010010010000: out_v[377] = 10'b0001101010;
    16'b0010000010110000: out_v[377] = 10'b1011001010;
    16'b0010010010110100: out_v[377] = 10'b0010011011;
    16'b0010011010100100: out_v[377] = 10'b0111001110;
    16'b0010010010010000: out_v[377] = 10'b1101011000;
    16'b0010111010100000: out_v[377] = 10'b0111111010;
    16'b0000010010000000: out_v[377] = 10'b0000101100;
    16'b0110010010000100: out_v[377] = 10'b0011011111;
    16'b0010011010100001: out_v[377] = 10'b0000001110;
    16'b0110110010110000: out_v[377] = 10'b0001011110;
    16'b0010010000000000: out_v[377] = 10'b0110011001;
    16'b0010000000100000: out_v[377] = 10'b0010101000;
    16'b0000010010000100: out_v[377] = 10'b0010011010;
    16'b0010011010100000: out_v[377] = 10'b1101011011;
    16'b0010110010100100: out_v[377] = 10'b1001001000;
    16'b0010010000100000: out_v[377] = 10'b0010110010;
    16'b0010101010100001: out_v[377] = 10'b1111001011;
    16'b0010010010110000: out_v[377] = 10'b0011011011;
    16'b0110010010100100: out_v[377] = 10'b1110010100;
    16'b0010000010100100: out_v[377] = 10'b0101101011;
    16'b0010000000110000: out_v[377] = 10'b1001101110;
    16'b0010110000100001: out_v[377] = 10'b0110111000;
    16'b0110010010100000: out_v[377] = 10'b1001000111;
    16'b0110010000100000: out_v[377] = 10'b0011100111;
    16'b0110010010000000: out_v[377] = 10'b0110111000;
    16'b0100101010100100: out_v[377] = 10'b0101111111;
    16'b0110010000110000: out_v[377] = 10'b0010011010;
    16'b0010101010100100: out_v[377] = 10'b1011011010;
    16'b0110011010100000: out_v[377] = 10'b1001000011;
    16'b0110000010000000: out_v[377] = 10'b1001000111;
    16'b0100111010100100: out_v[377] = 10'b0101011011;
    16'b0110000010100000: out_v[377] = 10'b1000111111;
    16'b0000101010100100: out_v[377] = 10'b1101011011;
    16'b0100010000110000: out_v[377] = 10'b0110011011;
    16'b0100101010100000: out_v[377] = 10'b1100001110;
    16'b0100010010100000: out_v[377] = 10'b1101000011;
    16'b0100010010110000: out_v[377] = 10'b1010001101;
    16'b0000101010100000: out_v[377] = 10'b1100001001;
    16'b0100011010100000: out_v[377] = 10'b0101011011;
    16'b0100011000100000: out_v[377] = 10'b0011010101;
    16'b0110101010100100: out_v[377] = 10'b1011010111;
    16'b0110101010100000: out_v[377] = 10'b0110011101;
    16'b0100001010100000: out_v[377] = 10'b0111010111;
    16'b0100000010100000: out_v[377] = 10'b1101111011;
    16'b0110010000000000: out_v[377] = 10'b0010010001;
    16'b0100111010100000: out_v[377] = 10'b0010110011;
    16'b0110010010110000: out_v[377] = 10'b1010011001;
    16'b0110000000000000: out_v[377] = 10'b0011010011;
    16'b0000101000100000: out_v[377] = 10'b0010000111;
    16'b0110000000100000: out_v[377] = 10'b0010101111;
    16'b0000010010110000: out_v[377] = 10'b0111010111;
    16'b0000011010100000: out_v[377] = 10'b0001011011;
    16'b0110100010100000: out_v[377] = 10'b1101100000;
    16'b0000000010100000: out_v[377] = 10'b0110011011;
    16'b0110111010100000: out_v[377] = 10'b0100111011;
    16'b0000010000110000: out_v[377] = 10'b1100010111;
    16'b0000000000100000: out_v[377] = 10'b1001011001;
    16'b0000010010100000: out_v[377] = 10'b0111010110;
    16'b0000011000100000: out_v[377] = 10'b0100011000;
    16'b0110111010100100: out_v[377] = 10'b1100010000;
    16'b0000101010000000: out_v[377] = 10'b0010100000;
    16'b0100011010010100: out_v[377] = 10'b1001110111;
    16'b0000001010000100: out_v[377] = 10'b1010111100;
    16'b0100111010000000: out_v[377] = 10'b1001100010;
    16'b0100110010010000: out_v[377] = 10'b1001111000;
    16'b0100011010000100: out_v[377] = 10'b0111000111;
    16'b0110000000110000: out_v[377] = 10'b0010110001;
    16'b0100010010000000: out_v[377] = 10'b1000001111;
    16'b0001101010000000: out_v[377] = 10'b1010001011;
    16'b0000011010000000: out_v[377] = 10'b0011100101;
    16'b0000011010000100: out_v[377] = 10'b0001100111;
    16'b0000001010000000: out_v[377] = 10'b1001110000;
    16'b0010101010000001: out_v[377] = 10'b1010110110;
    16'b0000111010000000: out_v[377] = 10'b0010110111;
    16'b0000101010000001: out_v[377] = 10'b1110001001;
    16'b0001111010000000: out_v[377] = 10'b1000100111;
    16'b0100010010010000: out_v[377] = 10'b0101110110;
    16'b0100010010000100: out_v[377] = 10'b0011110111;
    16'b0100110010000000: out_v[377] = 10'b0011110011;
    16'b0100111010000001: out_v[377] = 10'b1010011101;
    16'b0100001010000100: out_v[377] = 10'b1011101110;
    16'b0100011010000000: out_v[377] = 10'b0000111110;
    16'b0100011010010000: out_v[377] = 10'b0011100111;
    16'b0101011010000100: out_v[377] = 10'b1011011111;
    16'b0000100000000000: out_v[377] = 10'b0001000001;
    16'b0100110010100000: out_v[377] = 10'b0111001111;
    16'b0000100010100000: out_v[377] = 10'b1100011000;
    16'b0100100010000000: out_v[377] = 10'b1011010010;
    16'b0100100010100000: out_v[377] = 10'b0100101010;
    16'b0100110000010000: out_v[377] = 10'b1001000000;
    16'b0100100010010000: out_v[377] = 10'b1010111011;
    16'b0100100000100000: out_v[377] = 10'b0101011100;
    16'b0100100010110000: out_v[377] = 10'b1111110001;
    16'b0000110010010000: out_v[377] = 10'b1111111001;
    16'b0010100000100100: out_v[377] = 10'b1111100010;
    16'b0110011000100000: out_v[377] = 10'b1010101101;
    16'b0110111000100100: out_v[377] = 10'b0010101101;
    16'b0100101000100100: out_v[377] = 10'b1111001111;
    16'b0110100000100100: out_v[377] = 10'b0011100111;
    16'b0100000000100000: out_v[377] = 10'b1100101001;
    16'b0100100000100100: out_v[377] = 10'b0111110000;
    16'b0110010000100100: out_v[377] = 10'b1101110101;
    16'b0110110000100100: out_v[377] = 10'b0010110011;
    16'b0010101000100000: out_v[377] = 10'b1100010111;
    16'b0000100000100100: out_v[377] = 10'b0011111100;
    16'b0110100000100000: out_v[377] = 10'b1011111010;
    16'b0100111000100100: out_v[377] = 10'b1011011100;
    16'b0100101000100000: out_v[377] = 10'b0010110111;
    16'b0010101000100100: out_v[377] = 10'b0011101101;
    16'b0000101000100100: out_v[377] = 10'b0111000011;
    16'b0100010000100100: out_v[377] = 10'b0010111010;
    16'b0110101000100100: out_v[377] = 10'b1101000011;
    16'b0100110000100100: out_v[377] = 10'b0110010111;
    16'b0010100000000100: out_v[377] = 10'b0111111100;
    16'b0110101000100000: out_v[377] = 10'b1011000011;
    16'b0000110000100100: out_v[377] = 10'b1011111001;
    16'b0100001010100100: out_v[377] = 10'b0001011110;
    16'b0110100010000000: out_v[377] = 10'b1101111100;
    16'b0110001010100100: out_v[377] = 10'b1011110111;
    16'b0000001010100000: out_v[377] = 10'b0110010001;
    16'b0110111010110000: out_v[377] = 10'b0101101111;
    16'b0010001010000100: out_v[377] = 10'b1111001010;
    16'b0110000010110000: out_v[377] = 10'b0111000010;
    16'b0000101010100001: out_v[377] = 10'b0101011010;
    16'b0110100010100100: out_v[377] = 10'b1001111111;
    16'b0110001010100000: out_v[377] = 10'b0011100101;
    16'b0110110010010000: out_v[377] = 10'b0110001011;
    16'b0010001010100100: out_v[377] = 10'b0011011100;
    16'b0110010010010000: out_v[377] = 10'b0100001011;
    16'b0110011010100100: out_v[377] = 10'b0001011110;
    16'b0000000010100100: out_v[377] = 10'b1101101011;
    16'b0000001010100100: out_v[377] = 10'b0100010011;
    16'b0100000010100100: out_v[377] = 10'b0101001011;
    16'b0110110010100100: out_v[377] = 10'b1001111111;
    16'b0100100010100100: out_v[377] = 10'b1100001011;
    16'b0000100010100100: out_v[377] = 10'b1101001111;
    16'b0100010010100100: out_v[377] = 10'b1001011011;
    16'b0100110010100100: out_v[377] = 10'b0100011110;
    16'b0110000010100100: out_v[377] = 10'b1011110110;
    default: out_v[377] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000001000010: out_v[378] = 10'b1010111111;
    16'b0100100000000010: out_v[378] = 10'b0001001011;
    16'b0110100000000010: out_v[378] = 10'b0000110100;
    16'b0110000000010010: out_v[378] = 10'b1110100001;
    16'b0000000000000010: out_v[378] = 10'b1001001111;
    16'b0100000000000110: out_v[378] = 10'b1101000101;
    16'b0010000000000010: out_v[378] = 10'b1010100111;
    16'b0110000000000000: out_v[378] = 10'b0000011111;
    16'b0010100000010000: out_v[378] = 10'b0000010111;
    16'b0010000000000000: out_v[378] = 10'b0001110111;
    16'b0110000001000000: out_v[378] = 10'b0010000001;
    16'b0100000000000100: out_v[378] = 10'b1101010011;
    16'b0000100000010010: out_v[378] = 10'b0000010111;
    16'b0100100000010010: out_v[378] = 10'b0010001111;
    16'b0110000000000010: out_v[378] = 10'b0110100111;
    16'b0100000000000010: out_v[378] = 10'b1011000011;
    16'b0110000001000010: out_v[378] = 10'b1110000101;
    16'b0100000001000010: out_v[378] = 10'b1001011111;
    16'b0110000000000110: out_v[378] = 10'b1101000110;
    16'b0000000000000110: out_v[378] = 10'b0110010010;
    16'b0000000000010010: out_v[378] = 10'b1000111100;
    16'b0010100000000000: out_v[378] = 10'b1011001011;
    16'b0010000001000000: out_v[378] = 10'b0110100001;
    16'b0000100000000010: out_v[378] = 10'b0101010011;
    16'b0100100000010110: out_v[378] = 10'b0101001011;
    16'b0010100000010010: out_v[378] = 10'b1110001011;
    16'b0010100000000010: out_v[378] = 10'b1011110110;
    16'b0110100000010010: out_v[378] = 10'b1110110111;
    16'b0100000000010010: out_v[378] = 10'b0111110001;
    16'b0110100000000000: out_v[378] = 10'b1110100011;
    16'b0010000001000010: out_v[378] = 10'b1010110001;
    16'b0000100000010110: out_v[378] = 10'b0010010110;
    16'b0100100000000110: out_v[378] = 10'b1010001101;
    16'b0100000000010110: out_v[378] = 10'b1001111101;
    16'b0000000000000100: out_v[378] = 10'b1111011010;
    16'b0000100000010100: out_v[378] = 10'b1110000110;
    16'b0000000000000000: out_v[378] = 10'b0010111010;
    16'b0000000000010000: out_v[378] = 10'b0111110011;
    16'b0000000001000100: out_v[378] = 10'b0001000110;
    16'b0000000000010100: out_v[378] = 10'b0111100011;
    16'b0000100000010000: out_v[378] = 10'b1001011100;
    16'b0000100000000000: out_v[378] = 10'b0011101100;
    16'b0000100000000100: out_v[378] = 10'b0110110100;
    16'b0000000001000000: out_v[378] = 10'b0100100010;
    16'b0010000000000110: out_v[378] = 10'b0010111000;
    16'b0100100000000100: out_v[378] = 10'b0101110010;
    16'b0100000000010100: out_v[378] = 10'b1110111010;
    16'b0100000000000000: out_v[378] = 10'b0110110100;
    16'b0000000010000100: out_v[378] = 10'b0001111100;
    16'b0100000001000000: out_v[378] = 10'b0101000111;
    16'b0100000001000100: out_v[378] = 10'b1010000001;
    16'b0100000000010000: out_v[378] = 10'b1110100100;
    16'b0000000010000000: out_v[378] = 10'b0110000010;
    16'b0110000000000100: out_v[378] = 10'b0011001010;
    16'b0100000010000000: out_v[378] = 10'b0001010111;
    16'b0110000010000100: out_v[378] = 10'b1110000111;
    16'b0110000010000110: out_v[378] = 10'b1001000110;
    16'b0010000000000100: out_v[378] = 10'b1011011010;
    16'b0100100000010100: out_v[378] = 10'b0110011001;
    16'b0110000010000000: out_v[378] = 10'b0010001101;
    16'b0000000000010110: out_v[378] = 10'b1111101010;
    16'b0100000010000100: out_v[378] = 10'b0011100110;
    16'b0001000001000100: out_v[378] = 10'b0011110100;
    16'b0011000001000110: out_v[378] = 10'b0111011001;
    16'b0000000001000110: out_v[378] = 10'b1011101110;
    16'b0011000000000110: out_v[378] = 10'b1000001011;
    16'b0000100000000110: out_v[378] = 10'b0011111000;
    16'b0010000001000110: out_v[378] = 10'b0110011000;
    16'b0001000001000110: out_v[378] = 10'b1011011110;
    16'b0100000001000110: out_v[378] = 10'b1100011010;
    16'b0010100000000110: out_v[378] = 10'b0000111010;
    16'b0000100001000110: out_v[378] = 10'b0011111000;
    16'b0010100000000100: out_v[378] = 10'b1100111010;
    16'b0010100001000110: out_v[378] = 10'b1000100010;
    16'b0100100000000000: out_v[378] = 10'b1101010010;
    16'b0000100001000000: out_v[378] = 10'b1000100010;
    16'b0000100001000100: out_v[378] = 10'b0101101111;
    16'b0110000000010110: out_v[378] = 10'b0011010010;
    16'b0000001000000110: out_v[378] = 10'b1001011000;
    16'b0001000000000110: out_v[378] = 10'b0110110110;
    16'b0000001000000100: out_v[378] = 10'b1011001001;
    16'b0001000000000100: out_v[378] = 10'b1100110110;
    16'b0000101000000100: out_v[378] = 10'b0011101111;
    16'b0100100001000100: out_v[378] = 10'b0010100101;
    16'b0110000001000110: out_v[378] = 10'b1100011010;
    default: out_v[378] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000010000110: out_v[379] = 10'b0101110010;
    16'b0100001010000010: out_v[379] = 10'b1001100111;
    16'b0100000010100110: out_v[379] = 10'b0000101111;
    16'b0010000010000110: out_v[379] = 10'b1001001110;
    16'b0000000010100110: out_v[379] = 10'b0110110001;
    16'b0100000010100010: out_v[379] = 10'b0010100111;
    16'b0100000010100000: out_v[379] = 10'b1011000000;
    16'b0000000010000100: out_v[379] = 10'b0001001011;
    16'b0010000000000100: out_v[379] = 10'b0110110011;
    16'b0000000010100010: out_v[379] = 10'b1001001011;
    16'b0100000010000000: out_v[379] = 10'b1011110110;
    16'b0000000010100000: out_v[379] = 10'b0110101000;
    16'b0000001010000100: out_v[379] = 10'b0111010111;
    16'b0100000010000010: out_v[379] = 10'b0010011101;
    16'b0100000010000100: out_v[379] = 10'b1001100110;
    16'b0100000010000110: out_v[379] = 10'b1000011011;
    16'b0110000010000100: out_v[379] = 10'b1011011010;
    16'b0010000010100110: out_v[379] = 10'b1010110011;
    16'b0000000010100100: out_v[379] = 10'b0101001001;
    16'b0000001010100110: out_v[379] = 10'b0010101010;
    16'b0100000000100000: out_v[379] = 10'b0100001001;
    16'b0100000000100010: out_v[379] = 10'b0000000011;
    16'b0110000010000010: out_v[379] = 10'b1100110011;
    16'b0010000000000110: out_v[379] = 10'b1001110011;
    16'b0000010010000110: out_v[379] = 10'b0111011101;
    16'b0100000010100100: out_v[379] = 10'b0100011111;
    16'b0010000010000100: out_v[379] = 10'b1010110011;
    16'b0100001010100010: out_v[379] = 10'b0011001111;
    16'b0110000010100110: out_v[379] = 10'b1000010111;
    16'b0110000010000110: out_v[379] = 10'b1001100101;
    16'b0000000000000110: out_v[379] = 10'b1010100011;
    16'b0100000000000010: out_v[379] = 10'b0011011001;
    16'b0000000010000010: out_v[379] = 10'b0011111011;
    16'b0100001010100110: out_v[379] = 10'b1011100011;
    16'b0000010010100110: out_v[379] = 10'b1001011011;
    16'b0000001010100000: out_v[379] = 10'b0011111011;
    16'b0000000010000000: out_v[379] = 10'b1001100101;
    16'b0010000000100110: out_v[379] = 10'b1010011101;
    16'b0000001010100100: out_v[379] = 10'b1101000111;
    16'b0000000000000100: out_v[379] = 10'b0011001101;
    16'b0000100000100010: out_v[379] = 10'b1100110110;
    16'b0000100000100000: out_v[379] = 10'b0011100011;
    16'b0000100000000000: out_v[379] = 10'b0111001101;
    16'b0010100000000000: out_v[379] = 10'b0111100101;
    16'b0010100010000000: out_v[379] = 10'b0010010011;
    16'b0000100010000000: out_v[379] = 10'b1000011111;
    16'b0000101000100000: out_v[379] = 10'b0001110110;
    16'b0000000000100000: out_v[379] = 10'b1001101110;
    16'b0000100010100000: out_v[379] = 10'b1101100000;
    16'b0100100000100000: out_v[379] = 10'b0011000010;
    16'b0000101000100010: out_v[379] = 10'b1101001110;
    16'b0000100000000010: out_v[379] = 10'b1110001000;
    16'b0010100000100000: out_v[379] = 10'b1001001011;
    16'b0000000000000000: out_v[379] = 10'b1111000111;
    16'b0110100010000000: out_v[379] = 10'b0001101000;
    16'b0010000010000000: out_v[379] = 10'b1010011111;
    16'b0100100010000000: out_v[379] = 10'b1000100111;
    16'b0110100010100000: out_v[379] = 10'b0111110010;
    16'b0010100010100000: out_v[379] = 10'b0100011110;
    16'b0110100000000010: out_v[379] = 10'b1000100100;
    16'b0110100000100100: out_v[379] = 10'b0110001101;
    16'b0010100000100100: out_v[379] = 10'b1100001101;
    16'b0110100000000000: out_v[379] = 10'b1100011101;
    16'b0110100000100010: out_v[379] = 10'b1000100110;
    16'b0100100010100110: out_v[379] = 10'b1000101101;
    16'b0100100000000010: out_v[379] = 10'b1011100110;
    16'b0000100010100100: out_v[379] = 10'b0110001001;
    16'b0110000000100000: out_v[379] = 10'b1000001100;
    16'b0100100000010010: out_v[379] = 10'b0100011000;
    16'b0100100000100010: out_v[379] = 10'b1001001101;
    16'b0110000000000010: out_v[379] = 10'b1011101111;
    16'b0110100010000110: out_v[379] = 10'b0111100110;
    16'b0000100010100110: out_v[379] = 10'b0110001100;
    16'b0110100000100000: out_v[379] = 10'b1000001101;
    16'b0100100010000010: out_v[379] = 10'b0101011110;
    16'b0110000000000000: out_v[379] = 10'b1110011110;
    16'b0110000000100010: out_v[379] = 10'b1101011000;
    16'b0110100010100110: out_v[379] = 10'b1010010010;
    16'b0100100010100100: out_v[379] = 10'b1100001100;
    16'b0010100000100010: out_v[379] = 10'b1011111110;
    16'b0010100000000110: out_v[379] = 10'b0111001110;
    16'b0110000000000110: out_v[379] = 10'b0101110010;
    16'b0000100010000110: out_v[379] = 10'b1100001100;
    16'b0010100100000010: out_v[379] = 10'b1010001000;
    16'b0100100010000110: out_v[379] = 10'b0001001000;
    16'b0000100010000010: out_v[379] = 10'b1101100000;
    16'b0010100010100100: out_v[379] = 10'b0101001101;
    16'b0010100000000010: out_v[379] = 10'b1011011110;
    16'b0110100000010010: out_v[379] = 10'b0110001111;
    16'b0100100010000100: out_v[379] = 10'b0100100111;
    16'b0010000000100000: out_v[379] = 10'b0000011101;
    16'b0110100000000110: out_v[379] = 10'b0111111001;
    16'b0110000000010010: out_v[379] = 10'b1011110111;
    16'b0010100010000110: out_v[379] = 10'b0111100010;
    16'b0100100010100010: out_v[379] = 10'b1010100111;
    16'b0110100010100100: out_v[379] = 10'b1011011110;
    16'b0100100010010010: out_v[379] = 10'b1001001010;
    16'b0100101010100100: out_v[379] = 10'b0001011111;
    16'b0000101000100100: out_v[379] = 10'b1001011111;
    16'b0100100010100000: out_v[379] = 10'b0100111001;
    16'b0100110010100100: out_v[379] = 10'b0111100010;
    16'b0100100000100100: out_v[379] = 10'b1100011010;
    16'b0000110010100100: out_v[379] = 10'b1001011110;
    16'b0100101010100110: out_v[379] = 10'b0111101000;
    16'b0100101000100000: out_v[379] = 10'b0110000010;
    16'b0100101000000010: out_v[379] = 10'b1101011110;
    16'b0100101010000110: out_v[379] = 10'b0011011010;
    16'b0010000000100010: out_v[379] = 10'b1111011000;
    16'b0000101010000110: out_v[379] = 10'b1000111010;
    16'b0100101000100100: out_v[379] = 10'b1101010111;
    16'b0010000000000000: out_v[379] = 10'b1010111101;
    16'b0000101010100110: out_v[379] = 10'b1001011111;
    16'b0000101010100100: out_v[379] = 10'b1011001000;
    16'b0000100000100100: out_v[379] = 10'b0011010000;
    16'b0100101010000100: out_v[379] = 10'b0011110010;
    16'b0100100000000000: out_v[379] = 10'b1000111100;
    16'b0100110000000110: out_v[379] = 10'b0111110011;
    16'b0100110000100100: out_v[379] = 10'b0001011011;
    16'b0000100010000100: out_v[379] = 10'b1110111111;
    16'b0100101010000010: out_v[379] = 10'b1101010110;
    16'b0100000000000110: out_v[379] = 10'b1011000010;
    16'b0000101010000010: out_v[379] = 10'b0000010001;
    16'b0000100000000110: out_v[379] = 10'b1111011110;
    16'b0100100000000110: out_v[379] = 10'b1101001110;
    16'b0000100000000100: out_v[379] = 10'b1000100110;
    16'b0100110000100110: out_v[379] = 10'b1011101111;
    16'b0100110000100000: out_v[379] = 10'b1001110001;
    16'b0100010000000110: out_v[379] = 10'b1101101010;
    16'b0100110000000010: out_v[379] = 10'b1011101011;
    16'b0100100000000100: out_v[379] = 10'b1101110010;
    16'b0000101000000010: out_v[379] = 10'b1001011001;
    16'b0100010010000110: out_v[379] = 10'b0111001101;
    16'b0100100000100110: out_v[379] = 10'b0101010111;
    16'b0100000100000010: out_v[379] = 10'b0111011011;
    16'b0100110000100010: out_v[379] = 10'b1011110111;
    16'b0100110010000110: out_v[379] = 10'b1010001001;
    16'b0100010000000010: out_v[379] = 10'b0101010111;
    16'b0000100100000010: out_v[379] = 10'b0000111011;
    16'b0000101010000100: out_v[379] = 10'b0111001111;
    16'b0001000000100000: out_v[379] = 10'b1011111111;
    16'b0010100000000100: out_v[379] = 10'b0111100011;
    16'b0100101010100000: out_v[379] = 10'b1111111101;
    16'b0101100000100000: out_v[379] = 10'b0010000111;
    16'b0000110010000100: out_v[379] = 10'b0011011000;
    16'b0110100010000100: out_v[379] = 10'b0110110011;
    16'b0100101010000000: out_v[379] = 10'b0110100111;
    16'b0100110010000100: out_v[379] = 10'b1011000111;
    16'b0010100010000100: out_v[379] = 10'b0001000011;
    16'b0000000000000010: out_v[379] = 10'b1110110001;
    16'b0110100000000100: out_v[379] = 10'b1000100011;
    16'b0100001010000100: out_v[379] = 10'b1100100101;
    16'b0000000000100010: out_v[379] = 10'b1001010001;
    16'b0000100010010000: out_v[379] = 10'b0111111011;
    16'b0100000010010000: out_v[379] = 10'b1011111011;
    16'b0100100010010000: out_v[379] = 10'b0011011111;
    16'b0100000000000000: out_v[379] = 10'b1001010001;
    16'b0000000000010000: out_v[379] = 10'b1001011001;
    16'b0100000000110000: out_v[379] = 10'b1001100000;
    16'b0100100010010100: out_v[379] = 10'b0110110011;
    16'b0110000010000000: out_v[379] = 10'b1100110010;
    16'b0100100000110000: out_v[379] = 10'b0001101011;
    16'b0100000000010000: out_v[379] = 10'b1001000100;
    16'b0100100000010000: out_v[379] = 10'b0011101111;
    16'b0000100000010000: out_v[379] = 10'b0111000001;
    16'b0000000010010000: out_v[379] = 10'b1111010001;
    16'b0110100010000010: out_v[379] = 10'b1101100010;
    16'b0000100000110000: out_v[379] = 10'b0010011011;
    16'b0000100010010100: out_v[379] = 10'b0111000100;
    16'b0100101011100110: out_v[379] = 10'b0111001111;
    16'b0100000000100110: out_v[379] = 10'b0011110010;
    16'b0000101011100110: out_v[379] = 10'b0100110001;
    16'b0100001011100110: out_v[379] = 10'b0011110110;
    16'b0100010010100110: out_v[379] = 10'b0001011110;
    16'b0000101011100010: out_v[379] = 10'b0111011001;
    16'b0000100010100010: out_v[379] = 10'b0111100100;
    16'b0100110010100110: out_v[379] = 10'b0010100001;
    16'b0100000011100110: out_v[379] = 10'b0011111101;
    16'b0100010010100100: out_v[379] = 10'b0111011011;
    16'b0000101010100010: out_v[379] = 10'b1111001001;
    16'b0100010000100010: out_v[379] = 10'b0001111111;
    16'b0000100011100110: out_v[379] = 10'b0001110111;
    16'b0100100011100110: out_v[379] = 10'b0110010111;
    16'b0100101010100010: out_v[379] = 10'b1000000010;
    16'b0100110110100110: out_v[379] = 10'b1100001111;
    16'b0100110010100000: out_v[379] = 10'b1010000000;
    default: out_v[379] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1000001100101000: out_v[380] = 10'b1111110101;
    16'b1000001100111100: out_v[380] = 10'b0110110011;
    16'b1000001100000100: out_v[380] = 10'b1110011001;
    16'b1000000100111000: out_v[380] = 10'b0100011111;
    16'b1000001100111000: out_v[380] = 10'b1111101000;
    16'b0001001100011000: out_v[380] = 10'b1011111100;
    16'b0000011000100100: out_v[380] = 10'b1010010111;
    16'b1001001100111000: out_v[380] = 10'b0110101110;
    16'b1000001110101000: out_v[380] = 10'b1100111110;
    16'b1000001110001000: out_v[380] = 10'b1001011111;
    16'b1000001110000000: out_v[380] = 10'b1011010101;
    16'b1000001100011000: out_v[380] = 10'b0001000111;
    16'b1001001100111100: out_v[380] = 10'b1100100011;
    16'b1000001100101100: out_v[380] = 10'b1111101110;
    16'b1000001100011100: out_v[380] = 10'b0111101110;
    16'b0001001100111000: out_v[380] = 10'b0110111101;
    16'b1000001100001100: out_v[380] = 10'b1100111011;
    16'b1000001110011000: out_v[380] = 10'b0011011010;
    16'b1001001100011100: out_v[380] = 10'b1111001010;
    16'b0000001100101000: out_v[380] = 10'b1000101101;
    16'b1000001100100100: out_v[380] = 10'b0100000111;
    16'b1000001110111000: out_v[380] = 10'b1111101000;
    16'b1000001000101000: out_v[380] = 10'b1010001011;
    16'b1010001100101000: out_v[380] = 10'b1110010111;
    16'b0001001110011000: out_v[380] = 10'b0111101111;
    16'b0000001100101100: out_v[380] = 10'b1110011010;
    16'b1000001100001000: out_v[380] = 10'b1100100011;
    16'b0000011100101100: out_v[380] = 10'b0111010011;
    16'b1001001110011000: out_v[380] = 10'b0111110110;
    16'b1001001100011000: out_v[380] = 10'b0011111110;
    16'b1000001000111000: out_v[380] = 10'b1001111010;
    16'b1000000100101000: out_v[380] = 10'b0100101011;
    16'b1000011100111100: out_v[380] = 10'b1111111001;
    16'b0000001100100100: out_v[380] = 10'b1001011111;
    16'b1000011100101100: out_v[380] = 10'b0111010011;
    16'b1000001100000000: out_v[380] = 10'b0100001111;
    16'b0010011001000000: out_v[380] = 10'b0010100010;
    16'b0010011101000000: out_v[380] = 10'b1011000000;
    16'b0010000011100000: out_v[380] = 10'b0010011111;
    16'b0010000001100000: out_v[380] = 10'b0011110110;
    16'b0010001001100100: out_v[380] = 10'b0110010001;
    16'b0010001001000000: out_v[380] = 10'b1110011011;
    16'b0010001001000100: out_v[380] = 10'b1110010111;
    16'b0010000001000000: out_v[380] = 10'b0011001111;
    16'b0010000000100000: out_v[380] = 10'b1110010111;
    16'b0010010001000000: out_v[380] = 10'b1000100110;
    16'b0010010101000000: out_v[380] = 10'b0010111111;
    16'b0010001011100000: out_v[380] = 10'b0101001111;
    16'b0010011001100100: out_v[380] = 10'b0011100110;
    16'b0010001001100000: out_v[380] = 10'b0110100111;
    16'b0000000001100000: out_v[380] = 10'b1010001010;
    16'b0010011001000100: out_v[380] = 10'b0101000010;
    16'b0010001011000000: out_v[380] = 10'b1101010110;
    16'b0010011001100000: out_v[380] = 10'b1001100001;
    16'b0010011011100000: out_v[380] = 10'b1111101001;
    16'b0010011011000000: out_v[380] = 10'b0010011110;
    16'b0000001101101100: out_v[380] = 10'b1001001110;
    16'b0010011000100000: out_v[380] = 10'b1000100111;
    16'b0010011001001100: out_v[380] = 10'b1110110100;
    16'b0010011001101100: out_v[380] = 10'b1010101011;
    16'b0000011001100100: out_v[380] = 10'b0010001101;
    16'b0000011001100000: out_v[380] = 10'b0101001101;
    16'b0000011001101000: out_v[380] = 10'b0111100000;
    16'b0010011001101000: out_v[380] = 10'b0111010100;
    16'b0010011101101100: out_v[380] = 10'b1110010010;
    16'b0000011100100100: out_v[380] = 10'b1011010111;
    16'b1000001101101100: out_v[380] = 10'b1001110110;
    16'b1000001101101000: out_v[380] = 10'b1010100110;
    16'b0000010000100000: out_v[380] = 10'b1100111110;
    16'b0000011000101100: out_v[380] = 10'b0110010101;
    16'b0010011000100100: out_v[380] = 10'b0001110011;
    16'b0000011001101100: out_v[380] = 10'b1111001111;
    16'b0000011101101000: out_v[380] = 10'b0010110111;
    16'b0010001001101000: out_v[380] = 10'b1011101111;
    16'b0000011000100000: out_v[380] = 10'b1000010111;
    16'b0010011101101000: out_v[380] = 10'b1100011100;
    16'b0010011001001000: out_v[380] = 10'b0011000011;
    16'b0000011100100000: out_v[380] = 10'b0011110010;
    16'b0010011101100100: out_v[380] = 10'b1001110001;
    16'b0010001001101100: out_v[380] = 10'b1000110001;
    16'b0000011101001100: out_v[380] = 10'b1000001001;
    16'b0000011101101100: out_v[380] = 10'b1000111101;
    16'b0000011101001000: out_v[380] = 10'b0001101111;
    16'b0010010001100000: out_v[380] = 10'b1001001011;
    16'b0000000101101100: out_v[380] = 10'b1010111110;
    16'b0000011101000100: out_v[380] = 10'b1101110000;
    16'b0000011001001000: out_v[380] = 10'b0101111110;
    16'b0000010101101100: out_v[380] = 10'b1010110111;
    16'b0000011101100100: out_v[380] = 10'b0010101101;
    16'b0010011101100000: out_v[380] = 10'b0111001011;
    16'b0010011101000100: out_v[380] = 10'b0111001110;
    16'b0000011101100000: out_v[380] = 10'b1100011111;
    16'b0010011111000000: out_v[380] = 10'b0101010101;
    16'b0000001101101000: out_v[380] = 10'b1011100110;
    16'b0000010100101100: out_v[380] = 10'b1110011111;
    16'b0010011010000000: out_v[380] = 10'b0001100010;
    16'b0010011100000100: out_v[380] = 10'b1110111010;
    16'b0010010011000000: out_v[380] = 10'b1101101010;
    16'b0010011000000000: out_v[380] = 10'b1000100101;
    16'b0010001010000000: out_v[380] = 10'b0111011011;
    16'b0010001000100100: out_v[380] = 10'b1110011010;
    16'b0000001011000000: out_v[380] = 10'b0011110010;
    16'b0010011111100000: out_v[380] = 10'b0001011111;
    16'b0010011010100000: out_v[380] = 10'b1001100101;
    16'b0010011100100100: out_v[380] = 10'b0011111000;
    16'b0010001000000100: out_v[380] = 10'b0001011101;
    16'b0010011100100000: out_v[380] = 10'b1101001010;
    16'b0010010010000000: out_v[380] = 10'b0011011001;
    16'b0010010000000000: out_v[380] = 10'b1001011100;
    16'b0010011110000000: out_v[380] = 10'b0101011010;
    16'b0010011100101100: out_v[380] = 10'b1000001010;
    16'b0010001000000000: out_v[380] = 10'b1001110011;
    16'b0010011000000100: out_v[380] = 10'b1011000100;
    16'b0010001000100000: out_v[380] = 10'b0111011001;
    16'b0010011000001100: out_v[380] = 10'b0011001110;
    16'b0010011000101100: out_v[380] = 10'b0110110100;
    16'b0010000011000000: out_v[380] = 10'b0001010001;
    16'b0000010111110000: out_v[380] = 10'b0100011111;
    16'b0010011001110000: out_v[380] = 10'b0001011011;
    16'b0000010001010000: out_v[380] = 10'b1100010110;
    16'b0000010101011000: out_v[380] = 10'b1100111101;
    16'b0010010101100000: out_v[380] = 10'b1110001010;
    16'b0000010001100000: out_v[380] = 10'b1100011111;
    16'b0000010101001000: out_v[380] = 10'b0111010110;
    16'b0000010001000000: out_v[380] = 10'b1101010111;
    16'b0010010101010000: out_v[380] = 10'b1001011101;
    16'b0010010111100000: out_v[380] = 10'b1111011101;
    16'b0000010101101000: out_v[380] = 10'b1011010001;
    16'b0000010101100000: out_v[380] = 10'b0100110111;
    16'b0000010001101000: out_v[380] = 10'b0111010111;
    16'b0010010011100000: out_v[380] = 10'b0110110011;
    16'b0000010101110000: out_v[380] = 10'b1100100101;
    16'b1000010101111000: out_v[380] = 10'b1110101011;
    16'b0000000101010000: out_v[380] = 10'b1011111010;
    16'b0010011001010000: out_v[380] = 10'b0011110110;
    16'b0010010001010000: out_v[380] = 10'b1001100100;
    16'b0000010100101000: out_v[380] = 10'b1111011000;
    16'b0000010101000000: out_v[380] = 10'b1011010011;
    16'b0000011001010000: out_v[380] = 10'b0111010111;
    16'b0000010000000000: out_v[380] = 10'b0010010101;
    16'b0000010101111000: out_v[380] = 10'b1111001011;
    16'b1000000101011000: out_v[380] = 10'b0010011011;
    16'b0010010101110000: out_v[380] = 10'b1100110111;
    16'b0000010011100000: out_v[380] = 10'b1101011110;
    16'b0000011001000000: out_v[380] = 10'b1110001001;
    16'b0000010111100000: out_v[380] = 10'b0011111000;
    16'b0000010001110000: out_v[380] = 10'b1001111011;
    16'b0010010000100000: out_v[380] = 10'b1100011111;
    16'b0000010100111000: out_v[380] = 10'b0100111010;
    16'b0000010111111000: out_v[380] = 10'b1101110111;
    16'b0010010001101000: out_v[380] = 10'b1101001110;
    16'b0000010101010000: out_v[380] = 10'b1110011101;
    16'b0000010111101000: out_v[380] = 10'b1011010111;
    16'b0010011010010000: out_v[380] = 10'b0011011100;
    16'b0000000101100000: out_v[380] = 10'b1110100001;
    16'b0000001011100000: out_v[380] = 10'b1001101101;
    16'b0000001001000000: out_v[380] = 10'b1011100111;
    16'b0000001001100000: out_v[380] = 10'b1010110010;
    16'b0000000100100000: out_v[380] = 10'b0000110101;
    16'b0000001111100000: out_v[380] = 10'b0001100000;
    16'b0000001101100000: out_v[380] = 10'b1100110110;
    16'b0000001010000000: out_v[380] = 10'b0001011111;
    16'b0000000101101000: out_v[380] = 10'b1000101010;
    16'b0010000101101000: out_v[380] = 10'b1011111000;
    16'b0000001000100000: out_v[380] = 10'b1001111000;
    16'b0000000101000000: out_v[380] = 10'b0001100010;
    16'b0010000100100000: out_v[380] = 10'b0101101101;
    16'b0000001001100100: out_v[380] = 10'b0110111101;
    16'b0000000101110000: out_v[380] = 10'b0101100110;
    16'b0000001011010000: out_v[380] = 10'b0010110110;
    16'b0000000111100000: out_v[380] = 10'b1101110101;
    16'b0000001001000100: out_v[380] = 10'b1010111010;
    16'b0010010100100000: out_v[380] = 10'b0001111110;
    16'b0010000101100000: out_v[380] = 10'b0100100100;
    16'b1010011010010000: out_v[380] = 10'b0011110010;
    16'b0010010100101000: out_v[380] = 10'b0111100010;
    16'b0000001111000000: out_v[380] = 10'b0101011000;
    16'b0010011000101000: out_v[380] = 10'b1010100110;
    16'b0000001001101100: out_v[380] = 10'b0010110011;
    16'b0000001000101100: out_v[380] = 10'b1101000100;
    16'b1010010001100000: out_v[380] = 10'b0011001001;
    16'b1011010001111000: out_v[380] = 10'b1011101101;
    16'b1000011001101100: out_v[380] = 10'b0111101010;
    16'b0000001000000100: out_v[380] = 10'b0011000111;
    16'b0000001000100100: out_v[380] = 10'b1101001000;
    16'b0000000000100000: out_v[380] = 10'b1111001011;
    16'b1010011001101100: out_v[380] = 10'b1111000010;
    16'b1010010101111000: out_v[380] = 10'b0000111010;
    16'b0000001001101000: out_v[380] = 10'b0011001111;
    16'b0010010001100100: out_v[380] = 10'b1111000001;
    16'b1000010000100000: out_v[380] = 10'b0111000011;
    16'b1000010001100000: out_v[380] = 10'b0100110111;
    16'b0000000001000100: out_v[380] = 10'b1011111100;
    16'b1000001001101100: out_v[380] = 10'b1110111110;
    16'b1010011001100100: out_v[380] = 10'b1110011011;
    16'b1000000000100000: out_v[380] = 10'b0011100000;
    16'b1010010001101100: out_v[380] = 10'b1110011111;
    16'b0000000001100100: out_v[380] = 10'b1111011001;
    16'b1010010001111000: out_v[380] = 10'b1111101011;
    16'b1000001000101100: out_v[380] = 10'b0000011111;
    16'b0000000000100100: out_v[380] = 10'b1001011010;
    16'b1010011001111100: out_v[380] = 10'b1011001010;
    16'b1000011001100100: out_v[380] = 10'b1110111001;
    16'b1010010001100100: out_v[380] = 10'b1000111011;
    16'b1010010001101000: out_v[380] = 10'b1111000010;
    16'b1010010000100000: out_v[380] = 10'b1010001110;
    16'b0000010110100000: out_v[380] = 10'b0101001110;
    16'b0000010100100000: out_v[380] = 10'b0111011001;
    16'b0000010010100000: out_v[380] = 10'b0110001110;
    16'b0000000100000000: out_v[380] = 10'b0010100110;
    16'b0000010100110000: out_v[380] = 10'b0110111001;
    16'b0000010110110000: out_v[380] = 10'b0110100001;
    16'b0000011010100000: out_v[380] = 10'b0000010111;
    16'b0010010010100000: out_v[380] = 10'b1111010101;
    16'b0010010110100000: out_v[380] = 10'b0110001101;
    16'b1000000100100000: out_v[380] = 10'b0111001000;
    16'b0000010100000000: out_v[380] = 10'b0111001001;
    16'b0000000110100000: out_v[380] = 10'b0111101000;
    16'b1000000110110000: out_v[380] = 10'b0111011111;
    16'b1000010110100000: out_v[380] = 10'b1111100010;
    16'b0000000110110000: out_v[380] = 10'b0011111111;
    16'b0000011110100000: out_v[380] = 10'b0111100011;
    16'b1000000110100000: out_v[380] = 10'b0011110111;
    16'b1010010110100000: out_v[380] = 10'b0110111110;
    16'b0010011111001000: out_v[380] = 10'b0111010100;
    16'b0000011111000000: out_v[380] = 10'b0100011111;
    16'b0010011101001100: out_v[380] = 10'b0110011011;
    16'b0000011101000000: out_v[380] = 10'b1111001010;
    16'b0000011111100000: out_v[380] = 10'b1111000001;
    16'b0000011011100000: out_v[380] = 10'b1101001011;
    16'b0010011101001000: out_v[380] = 10'b1110000001;
    16'b0010011111101000: out_v[380] = 10'b1001011000;
    16'b0000011011000000: out_v[380] = 10'b0110000010;
    16'b0010011111010000: out_v[380] = 10'b0110010110;
    16'b0010011110100000: out_v[380] = 10'b1001101011;
    16'b0010011111110000: out_v[380] = 10'b1001001010;
    16'b0000011111111000: out_v[380] = 10'b1001110111;
    16'b0000011111110000: out_v[380] = 10'b1101001011;
    16'b0010010111110000: out_v[380] = 10'b1111000100;
    16'b0010010001110000: out_v[380] = 10'b1100001010;
    16'b0000011101110000: out_v[380] = 10'b0011010010;
    default: out_v[380] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000001000010000: out_v[381] = 10'b0010100011;
    16'b0010001000000100: out_v[381] = 10'b1100010001;
    16'b0010001000000110: out_v[381] = 10'b0101011110;
    16'b0000001000000100: out_v[381] = 10'b1100010110;
    16'b0010001000010100: out_v[381] = 10'b1110010011;
    16'b0010000000000110: out_v[381] = 10'b1011111001;
    16'b0010000000000100: out_v[381] = 10'b0011100001;
    16'b0010000000000000: out_v[381] = 10'b0101100000;
    16'b0000001000010100: out_v[381] = 10'b0010010010;
    16'b0010001000000000: out_v[381] = 10'b1101000101;
    16'b0000001000000000: out_v[381] = 10'b0100011110;
    16'b0010001000010110: out_v[381] = 10'b1110010011;
    16'b0010001000010000: out_v[381] = 10'b0000111000;
    16'b0000001000000110: out_v[381] = 10'b0010111100;
    16'b0010000000000010: out_v[381] = 10'b0111100101;
    16'b0000000000010000: out_v[381] = 10'b0100001011;
    16'b0000001000010110: out_v[381] = 10'b1000011101;
    16'b1010001100000100: out_v[381] = 10'b1100001101;
    16'b0010000000010000: out_v[381] = 10'b0110010111;
    16'b0000000000000110: out_v[381] = 10'b0110111011;
    16'b0000000000000100: out_v[381] = 10'b0011110111;
    16'b0010000000010110: out_v[381] = 10'b0011001000;
    16'b0000000000000000: out_v[381] = 10'b0101101110;
    16'b1000000100000000: out_v[381] = 10'b1010110011;
    16'b0000000000000010: out_v[381] = 10'b1001011101;
    16'b1010001100000000: out_v[381] = 10'b1000011100;
    16'b0000000000010010: out_v[381] = 10'b1000101111;
    16'b1010000100010010: out_v[381] = 10'b0011000110;
    16'b0000001000010010: out_v[381] = 10'b0010100000;
    16'b1010001100010000: out_v[381] = 10'b1001111100;
    16'b1010000100010000: out_v[381] = 10'b1110110000;
    16'b0010001000010010: out_v[381] = 10'b1110011000;
    16'b0010001000000010: out_v[381] = 10'b0011111110;
    16'b0010000000010010: out_v[381] = 10'b0110001110;
    16'b1010001100000010: out_v[381] = 10'b0000100100;
    16'b1010000100000000: out_v[381] = 10'b0100011110;
    16'b1010000100000010: out_v[381] = 10'b1010010111;
    16'b1010001100010010: out_v[381] = 10'b1110011011;
    16'b0000001000000010: out_v[381] = 10'b0101011111;
    16'b1000000100000010: out_v[381] = 10'b1001100011;
    16'b0010000000010100: out_v[381] = 10'b1100110010;
    16'b0000000000010110: out_v[381] = 10'b0110000010;
    16'b0000000000010100: out_v[381] = 10'b1100100010;
    16'b0000000010000100: out_v[381] = 10'b1111100110;
    16'b1000001100000000: out_v[381] = 10'b1101000100;
    16'b1000001100000110: out_v[381] = 10'b0110010010;
    16'b1000001100010000: out_v[381] = 10'b1001100110;
    16'b1010001100010100: out_v[381] = 10'b1011001010;
    16'b1010000100000100: out_v[381] = 10'b1111101101;
    16'b1000001100000100: out_v[381] = 10'b1111111110;
    16'b0010011000010100: out_v[381] = 10'b1110001011;
    16'b0000010000010100: out_v[381] = 10'b1110011111;
    16'b1000000100000100: out_v[381] = 10'b1110001011;
    16'b1010000100010100: out_v[381] = 10'b1001011100;
    16'b1010001100000110: out_v[381] = 10'b1001001000;
    16'b1000000100000110: out_v[381] = 10'b0110100011;
    16'b1000001100010100: out_v[381] = 10'b0011010111;
    16'b1000001100000010: out_v[381] = 10'b1010110000;
    16'b0000010000010110: out_v[381] = 10'b0100000011;
    16'b1000000100010110: out_v[381] = 10'b1011001010;
    16'b0000011000010100: out_v[381] = 10'b1110101100;
    16'b1010000100010110: out_v[381] = 10'b1001110110;
    16'b1000000100010100: out_v[381] = 10'b0110011111;
    16'b0000001000000001: out_v[381] = 10'b1101111101;
    16'b0000000001010000: out_v[381] = 10'b1000001101;
    16'b0000000001000000: out_v[381] = 10'b1010101000;
    16'b0000000010010000: out_v[381] = 10'b1001001111;
    16'b0000001000010001: out_v[381] = 10'b0010110011;
    16'b0000000001010100: out_v[381] = 10'b0001100101;
    16'b0000001001010000: out_v[381] = 10'b0111111001;
    16'b0000001010000000: out_v[381] = 10'b0011001000;
    16'b0000000010010100: out_v[381] = 10'b1100101111;
    16'b0000001001010100: out_v[381] = 10'b1111010011;
    16'b0000000010000000: out_v[381] = 10'b0011011100;
    16'b0000001000010101: out_v[381] = 10'b1010100011;
    16'b0000001001000100: out_v[381] = 10'b1101111110;
    16'b0000001001000000: out_v[381] = 10'b1111100011;
    16'b0000001010010000: out_v[381] = 10'b0111111001;
    16'b0000000001000100: out_v[381] = 10'b0101111110;
    default: out_v[381] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000010010100000: out_v[382] = 10'b1001011111;
    16'b0100010011100000: out_v[382] = 10'b1001000101;
    16'b0100010001000000: out_v[382] = 10'b0100011011;
    16'b0100010000100000: out_v[382] = 10'b1010100111;
    16'b0100000011100000: out_v[382] = 10'b1101000110;
    16'b0100010010100000: out_v[382] = 10'b0010011011;
    16'b0000000011000000: out_v[382] = 10'b0110100011;
    16'b0100000001100000: out_v[382] = 10'b1110010001;
    16'b0100000001000000: out_v[382] = 10'b1001110111;
    16'b0100000010100000: out_v[382] = 10'b0010101100;
    16'b0000010011100000: out_v[382] = 10'b0010011111;
    16'b0000000011100000: out_v[382] = 10'b1100011100;
    16'b0000010000100000: out_v[382] = 10'b1100011000;
    16'b0000010010000000: out_v[382] = 10'b1001101111;
    16'b0000010011000000: out_v[382] = 10'b0100110111;
    16'b0100010000000000: out_v[382] = 10'b1001000110;
    16'b0100010010000000: out_v[382] = 10'b0000000101;
    16'b0100010001100000: out_v[382] = 10'b1100110011;
    16'b0100000011000000: out_v[382] = 10'b1001101101;
    16'b0100010011000000: out_v[382] = 10'b0011110101;
    16'b0000000010100000: out_v[382] = 10'b1101010001;
    16'b0100000011110000: out_v[382] = 10'b1010101110;
    16'b0000000011101100: out_v[382] = 10'b0011100101;
    16'b0100000001101100: out_v[382] = 10'b0100111101;
    16'b0100000001110000: out_v[382] = 10'b1100011011;
    16'b0100000000000000: out_v[382] = 10'b0011011100;
    16'b0000010000000000: out_v[382] = 10'b0010100001;
    16'b0000000010000000: out_v[382] = 10'b0110000111;
    16'b0000000011001100: out_v[382] = 10'b0101000111;
    16'b0100010001101100: out_v[382] = 10'b0011100001;
    16'b0000000000100000: out_v[382] = 10'b1000001010;
    16'b0100000000100000: out_v[382] = 10'b1011010011;
    16'b0100010010100010: out_v[382] = 10'b0110110010;
    16'b0000000000000000: out_v[382] = 10'b0010010111;
    16'b0000000000101100: out_v[382] = 10'b1000101101;
    16'b0000000000001100: out_v[382] = 10'b0011101010;
    16'b0100000010000000: out_v[382] = 10'b1001001110;
    16'b0000000000101000: out_v[382] = 10'b1011101101;
    16'b0100000000110000: out_v[382] = 10'b1111000101;
    16'b0100010010010000: out_v[382] = 10'b0110001011;
    16'b0100000010110000: out_v[382] = 10'b0111000011;
    16'b0100010000110000: out_v[382] = 10'b1100111110;
    16'b0100010010110000: out_v[382] = 10'b0111100111;
    16'b0100010010000010: out_v[382] = 10'b0101101110;
    16'b0100000010010000: out_v[382] = 10'b1110011011;
    16'b0100010011110000: out_v[382] = 10'b0000010101;
    16'b0100010001110000: out_v[382] = 10'b1001110110;
    16'b0100110000100000: out_v[382] = 10'b0010011001;
    16'b0100000010000010: out_v[382] = 10'b1111100111;
    16'b0100100000100000: out_v[382] = 10'b0001100111;
    16'b0100100000110000: out_v[382] = 10'b0010100111;
    16'b0100010011010000: out_v[382] = 10'b1011100011;
    16'b0000010001101100: out_v[382] = 10'b1011100101;
    16'b0000110000101100: out_v[382] = 10'b0010100110;
    16'b0100010000101100: out_v[382] = 10'b1100010011;
    16'b0000010000101000: out_v[382] = 10'b0100000111;
    16'b0000010000101100: out_v[382] = 10'b0011100010;
    16'b0000010000100010: out_v[382] = 10'b1100011011;
    16'b0000000001101100: out_v[382] = 10'b0110111000;
    16'b0000010001100000: out_v[382] = 10'b1011001000;
    16'b0000010000000010: out_v[382] = 10'b0001110100;
    16'b0000110000100000: out_v[382] = 10'b0111110110;
    16'b0000010010101100: out_v[382] = 10'b1110111110;
    16'b0100010000100010: out_v[382] = 10'b1101001101;
    16'b0000010001000000: out_v[382] = 10'b1110110000;
    16'b0000000001100000: out_v[382] = 10'b1001101010;
    16'b0000100000101100: out_v[382] = 10'b0100110101;
    16'b0000010001001100: out_v[382] = 10'b0010011111;
    16'b0000000001000000: out_v[382] = 10'b1010110000;
    16'b0000000001001100: out_v[382] = 10'b1111000001;
    16'b0000010000001100: out_v[382] = 10'b1100011000;
    16'b0000110000000000: out_v[382] = 10'b0001011010;
    16'b0000010011101100: out_v[382] = 10'b0011110011;
    16'b0100010001010000: out_v[382] = 10'b1001110010;
    16'b0100000001010000: out_v[382] = 10'b0011000000;
    16'b0110010010100000: out_v[382] = 10'b0101000010;
    16'b0000110001001100: out_v[382] = 10'b1000010111;
    16'b0000110001101100: out_v[382] = 10'b0011001001;
    16'b0000100001101100: out_v[382] = 10'b1111010001;
    16'b0000100001100000: out_v[382] = 10'b0001111011;
    16'b0100110001100000: out_v[382] = 10'b0111111010;
    16'b0000110001100000: out_v[382] = 10'b0111000000;
    16'b0000010001101000: out_v[382] = 10'b1011001110;
    16'b0100000000101100: out_v[382] = 10'b0101010100;
    16'b0100010001001100: out_v[382] = 10'b0110010010;
    16'b0100000001101000: out_v[382] = 10'b1111100100;
    16'b0100000001001100: out_v[382] = 10'b0110101111;
    16'b0100000000001100: out_v[382] = 10'b1100000110;
    16'b0100010000001100: out_v[382] = 10'b1111101000;
    default: out_v[382] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000000001000110: out_v[383] = 10'b0011100011;
    16'b0000000000000110: out_v[383] = 10'b1110101000;
    16'b0000000101000110: out_v[383] = 10'b0010100011;
    16'b0010000001000100: out_v[383] = 10'b1000000011;
    16'b0000000001000010: out_v[383] = 10'b0000111101;
    16'b0000000000000100: out_v[383] = 10'b1100100010;
    16'b0010000101000100: out_v[383] = 10'b1100000101;
    16'b0010000100000100: out_v[383] = 10'b0111000101;
    16'b0000000001000100: out_v[383] = 10'b0110000100;
    16'b0010000001000110: out_v[383] = 10'b1000001111;
    16'b0000000100000110: out_v[383] = 10'b0000111001;
    16'b0000000101000100: out_v[383] = 10'b0100001101;
    16'b0010000111000100: out_v[383] = 10'b0010001101;
    16'b0010000010000100: out_v[383] = 10'b1011001011;
    16'b0010000000000100: out_v[383] = 10'b0111001011;
    16'b0000000000000010: out_v[383] = 10'b0011010011;
    16'b0010000001000000: out_v[383] = 10'b1001001001;
    16'b0010000011000100: out_v[383] = 10'b1100100001;
    16'b0000000101000010: out_v[383] = 10'b1001001000;
    16'b0010000101000110: out_v[383] = 10'b0001100110;
    16'b0000000100000100: out_v[383] = 10'b0111001001;
    16'b0000000001000000: out_v[383] = 10'b0110110011;
    16'b0000000000000000: out_v[383] = 10'b0000011010;
    16'b0000000100000000: out_v[383] = 10'b0110011001;
    16'b0000000111000100: out_v[383] = 10'b0010010101;
    16'b0010000101000010: out_v[383] = 10'b1111100111;
    16'b0000000101000000: out_v[383] = 10'b1101000011;
    16'b0010000100000110: out_v[383] = 10'b1011100100;
    16'b0010000111000010: out_v[383] = 10'b0011000111;
    16'b0010000111000110: out_v[383] = 10'b0100000010;
    16'b0000000011000100: out_v[383] = 10'b1001110110;
    16'b0000000111000110: out_v[383] = 10'b1110100010;
    16'b0010000101000000: out_v[383] = 10'b0011001110;
    16'b0010000011000110: out_v[383] = 10'b0100000110;
    16'b0010000110000110: out_v[383] = 10'b0110100001;
    16'b0010000111000000: out_v[383] = 10'b1111100010;
    16'b0010000000000110: out_v[383] = 10'b0100100110;
    16'b0010000001000010: out_v[383] = 10'b0100000101;
    16'b0010000010000110: out_v[383] = 10'b0100101010;
    16'b0000000100000010: out_v[383] = 10'b0110111000;
    16'b0010000010000010: out_v[383] = 10'b1000111010;
    16'b0010000010000000: out_v[383] = 10'b1010011010;
    16'b0000000010000010: out_v[383] = 10'b0000011010;
    16'b0000000000010010: out_v[383] = 10'b1101110001;
    16'b0000000000010000: out_v[383] = 10'b1111001101;
    16'b0000010000000010: out_v[383] = 10'b1010000010;
    16'b0000000001010000: out_v[383] = 10'b0011011010;
    16'b0000000001010010: out_v[383] = 10'b0011111000;
    16'b0000000010000110: out_v[383] = 10'b0100010100;
    default: out_v[383] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0010100111101010: out_v[384] = 10'b1010011001;
    16'b0000100101101010: out_v[384] = 10'b0101100011;
    16'b1010100111000010: out_v[384] = 10'b1100100110;
    16'b1010100100000010: out_v[384] = 10'b1000010101;
    16'b0000000101101000: out_v[384] = 10'b1000001001;
    16'b0010100100000010: out_v[384] = 10'b0111001110;
    16'b0010100111001010: out_v[384] = 10'b1010011011;
    16'b0010100011101010: out_v[384] = 10'b1000100011;
    16'b0010100111000010: out_v[384] = 10'b0111110001;
    16'b0010100011000010: out_v[384] = 10'b1010101010;
    16'b1010100111101010: out_v[384] = 10'b0110010101;
    16'b0010100110000010: out_v[384] = 10'b1101000111;
    16'b1010000111000010: out_v[384] = 10'b1101001110;
    16'b1000000110000000: out_v[384] = 10'b1011011111;
    16'b1010000110000000: out_v[384] = 10'b1100000001;
    16'b0000100101101000: out_v[384] = 10'b1100111111;
    16'b0000000100101000: out_v[384] = 10'b0010010011;
    16'b0000100100101010: out_v[384] = 10'b1000011001;
    16'b1010100011000010: out_v[384] = 10'b0101011100;
    16'b0010100101101010: out_v[384] = 10'b0010110110;
    16'b1010100111100010: out_v[384] = 10'b0110001111;
    16'b1010100110000010: out_v[384] = 10'b1101110010;
    16'b1000000110000010: out_v[384] = 10'b1010010110;
    16'b1010000010000010: out_v[384] = 10'b1011001111;
    16'b0010100101100010: out_v[384] = 10'b0100011000;
    16'b1010100111001010: out_v[384] = 10'b1110000111;
    16'b1010000110000010: out_v[384] = 10'b0111010000;
    16'b1010100110100010: out_v[384] = 10'b1011111111;
    16'b1010100101101010: out_v[384] = 10'b0010101010;
    16'b0010100101000010: out_v[384] = 10'b0111100100;
    16'b1010100110101010: out_v[384] = 10'b1001111110;
    16'b1010100010000010: out_v[384] = 10'b1001001011;
    16'b0010100111101000: out_v[384] = 10'b1111101110;
    16'b0010100101101000: out_v[384] = 10'b1001011010;
    16'b1000100110000010: out_v[384] = 10'b0010101111;
    16'b0010100111100010: out_v[384] = 10'b1001100110;
    16'b0000000100101100: out_v[384] = 10'b0111100011;
    16'b0000010100000100: out_v[384] = 10'b1101110011;
    16'b0000010000000100: out_v[384] = 10'b1100100001;
    16'b0000010010000000: out_v[384] = 10'b1001100111;
    16'b0000010000000000: out_v[384] = 10'b1000111011;
    16'b0000010100000000: out_v[384] = 10'b1000111001;
    16'b0000010010100000: out_v[384] = 10'b1110100011;
    16'b0000010010100100: out_v[384] = 10'b0011101111;
    16'b0000010010000100: out_v[384] = 10'b1010100111;
    16'b0010010010000100: out_v[384] = 10'b0001110110;
    16'b0000010100100100: out_v[384] = 10'b1010001110;
    16'b0000010100001100: out_v[384] = 10'b0000011110;
    16'b0000010100101100: out_v[384] = 10'b1101000110;
    16'b0010010010100100: out_v[384] = 10'b1101000011;
    16'b0010010010100000: out_v[384] = 10'b1001110010;
    16'b0000010000100000: out_v[384] = 10'b1110001110;
    16'b0000010110000100: out_v[384] = 10'b0010110101;
    16'b1010110110000110: out_v[384] = 10'b0000110100;
    16'b1000010110000100: out_v[384] = 10'b0101010011;
    16'b1000110110000110: out_v[384] = 10'b0100001001;
    16'b1010010110000100: out_v[384] = 10'b1001110110;
    16'b1000010110000110: out_v[384] = 10'b1111011000;
    16'b1010110010000110: out_v[384] = 10'b1010001110;
    16'b0000110100000110: out_v[384] = 10'b0010110101;
    16'b0000110110000110: out_v[384] = 10'b1111101011;
    16'b0000010101000100: out_v[384] = 10'b0000010101;
    16'b1010110110001110: out_v[384] = 10'b0010001110;
    16'b1000110100000110: out_v[384] = 10'b0111110000;
    16'b0010110110000110: out_v[384] = 10'b1001001010;
    16'b0010010110000100: out_v[384] = 10'b0010111101;
    16'b1010100110000110: out_v[384] = 10'b0110011011;
    16'b1000110110001110: out_v[384] = 10'b0100011110;
    16'b1000110110000010: out_v[384] = 10'b0110111011;
    16'b0000110010000110: out_v[384] = 10'b1100001101;
    16'b1010010110000110: out_v[384] = 10'b0001011100;
    16'b1000100110000110: out_v[384] = 10'b1011100010;
    16'b1000110010000110: out_v[384] = 10'b0100101111;
    16'b1000110010000010: out_v[384] = 10'b0111111100;
    16'b0010010111000100: out_v[384] = 10'b0011111001;
    16'b1010110010000010: out_v[384] = 10'b0110101011;
    16'b0010100111001110: out_v[384] = 10'b1100110000;
    16'b0000110110001010: out_v[384] = 10'b0110001011;
    16'b0010110110001110: out_v[384] = 10'b0111001000;
    16'b1010110111101110: out_v[384] = 10'b0011101000;
    16'b0000100110101110: out_v[384] = 10'b0011001111;
    16'b1000100110101110: out_v[384] = 10'b1011011101;
    16'b0000010110001100: out_v[384] = 10'b1111001001;
    16'b1000100111101110: out_v[384] = 10'b1111010110;
    16'b0000110110001110: out_v[384] = 10'b1111100101;
    16'b1000110110101110: out_v[384] = 10'b1111010111;
    16'b0000100110001110: out_v[384] = 10'b1110000011;
    16'b0010110111001110: out_v[384] = 10'b1110000011;
    16'b0010010110001100: out_v[384] = 10'b1001000010;
    16'b1010110110101110: out_v[384] = 10'b0110110101;
    16'b0000100110101100: out_v[384] = 10'b0110011111;
    16'b0010100110001110: out_v[384] = 10'b0111011110;
    16'b0000100010101110: out_v[384] = 10'b1101011010;
    16'b1000110111001110: out_v[384] = 10'b1011110000;
    16'b1010010111001110: out_v[384] = 10'b0100110011;
    16'b1000110111101110: out_v[384] = 10'b1111101010;
    16'b0010100110101110: out_v[384] = 10'b0110011110;
    16'b1000000011101110: out_v[384] = 10'b1010100111;
    16'b0010110110000100: out_v[384] = 10'b1011001001;
    16'b0010110110001100: out_v[384] = 10'b1111010001;
    16'b1000000111101110: out_v[384] = 10'b1111011111;
    16'b1010110111001110: out_v[384] = 10'b1010011000;
    16'b0010110110101110: out_v[384] = 10'b0110110000;
    16'b0010100111101110: out_v[384] = 10'b1001001011;
    16'b1010100111101110: out_v[384] = 10'b0110111011;
    16'b0000110110101110: out_v[384] = 10'b1110110000;
    16'b0000100111101110: out_v[384] = 10'b1011011110;
    16'b0000110100001100: out_v[384] = 10'b0001110111;
    16'b0010010100000100: out_v[384] = 10'b0010011001;
    16'b0010010010001100: out_v[384] = 10'b0111110011;
    16'b0000010000101000: out_v[384] = 10'b0000110010;
    16'b0010010101001100: out_v[384] = 10'b0011101111;
    16'b0010010000101100: out_v[384] = 10'b0011011101;
    16'b0000010101001100: out_v[384] = 10'b1100010010;
    16'b0010010011101100: out_v[384] = 10'b1001111101;
    16'b0010010000000100: out_v[384] = 10'b1010111000;
    16'b0010010000001100: out_v[384] = 10'b0111001011;
    16'b0010010110101100: out_v[384] = 10'b0101110000;
    16'b0010010000000000: out_v[384] = 10'b1001101110;
    16'b0000110100000100: out_v[384] = 10'b0011110101;
    16'b0010010001000100: out_v[384] = 10'b1101000101;
    16'b0010010100101100: out_v[384] = 10'b1111000010;
    16'b0000010000101100: out_v[384] = 10'b0001011001;
    16'b0000010101101100: out_v[384] = 10'b0001110100;
    16'b0010010100001100: out_v[384] = 10'b1011000011;
    16'b0010010101000100: out_v[384] = 10'b0111100011;
    16'b0000010000001100: out_v[384] = 10'b1110011001;
    16'b0010010101101100: out_v[384] = 10'b0010110110;
    16'b0000010001101100: out_v[384] = 10'b0011001010;
    16'b0010010111101100: out_v[384] = 10'b0100011011;
    16'b0010010001101100: out_v[384] = 10'b1011100101;
    16'b0010010010101100: out_v[384] = 10'b0001100111;
    16'b0010010111001100: out_v[384] = 10'b0110100111;
    16'b1000110100001110: out_v[384] = 10'b0010000101;
    16'b0010010010000000: out_v[384] = 10'b1010110110;
    16'b0000010010101100: out_v[384] = 10'b1101111011;
    16'b0010010011001100: out_v[384] = 10'b0110100011;
    16'b0000110100001110: out_v[384] = 10'b1110011111;
    16'b1000110101001110: out_v[384] = 10'b0001110011;
    16'b0010010011000100: out_v[384] = 10'b0111001010;
    16'b0000010001001100: out_v[384] = 10'b1101000110;
    16'b0000010100101000: out_v[384] = 10'b1101100000;
    16'b0010110110101010: out_v[384] = 10'b1010100011;
    16'b0000110100101000: out_v[384] = 10'b1110101101;
    16'b0010110100101010: out_v[384] = 10'b1100101011;
    16'b1010000011101110: out_v[384] = 10'b1011110010;
    16'b0010010100001000: out_v[384] = 10'b0101101011;
    16'b1010110010001010: out_v[384] = 10'b0001011101;
    16'b0010110010101110: out_v[384] = 10'b1101110001;
    16'b0010100010001110: out_v[384] = 10'b0100111111;
    16'b1010000011001110: out_v[384] = 10'b0001100110;
    16'b0000110100101010: out_v[384] = 10'b1101000110;
    16'b1010100011101110: out_v[384] = 10'b0000011011;
    16'b0000000000101000: out_v[384] = 10'b0011111100;
    16'b0010100011101110: out_v[384] = 10'b1111110010;
    16'b0000010100001000: out_v[384] = 10'b0111110100;
    16'b1010110110001010: out_v[384] = 10'b0011100000;
    16'b0010010100101000: out_v[384] = 10'b1110111100;
    16'b0010010110101000: out_v[384] = 10'b0110011000;
    16'b0010100010101110: out_v[384] = 10'b0011110101;
    16'b0010100110101100: out_v[384] = 10'b1001100110;
    16'b0000010100100000: out_v[384] = 10'b0110100100;
    16'b0010110110001010: out_v[384] = 10'b0001100110;
    16'b1010110110101010: out_v[384] = 10'b1111010000;
    16'b0000110000101010: out_v[384] = 10'b0111011111;
    16'b0000100000101010: out_v[384] = 10'b0111010100;
    16'b0000110011101110: out_v[384] = 10'b0111110011;
    16'b0010110010000110: out_v[384] = 10'b1001111010;
    16'b0010110011101110: out_v[384] = 10'b1010111111;
    16'b1010110011000010: out_v[384] = 10'b1110111000;
    16'b1010110011001110: out_v[384] = 10'b0100110111;
    16'b0000110000101110: out_v[384] = 10'b1001110111;
    16'b0000100001101010: out_v[384] = 10'b1011100111;
    16'b0000110101101110: out_v[384] = 10'b1101000011;
    16'b1010110011101110: out_v[384] = 10'b1001001000;
    16'b1010110011000110: out_v[384] = 10'b0011001011;
    16'b0010110001101110: out_v[384] = 10'b0110111111;
    16'b0000110001101110: out_v[384] = 10'b1110100101;
    16'b0010110011000110: out_v[384] = 10'b0001101110;
    16'b0010110011001110: out_v[384] = 10'b1011010010;
    16'b1010110010001110: out_v[384] = 10'b0110011111;
    16'b0000110100101110: out_v[384] = 10'b0101010000;
    16'b0000110101101010: out_v[384] = 10'b0011000011;
    16'b0000110001101010: out_v[384] = 10'b0110110111;
    16'b1000110000000110: out_v[384] = 10'b0101100000;
    16'b0000110000101000: out_v[384] = 10'b1101011111;
    16'b0000110001101100: out_v[384] = 10'b1110011111;
    16'b0000110000101100: out_v[384] = 10'b0010110101;
    16'b1010100011101010: out_v[384] = 10'b0100110111;
    16'b0010110010001110: out_v[384] = 10'b1111001001;
    16'b0000000100000000: out_v[384] = 10'b0010110111;
    16'b0010000110000100: out_v[384] = 10'b0100000101;
    16'b0010000100000100: out_v[384] = 10'b0101010101;
    16'b0000000100000100: out_v[384] = 10'b1000101111;
    16'b0010000100100100: out_v[384] = 10'b0111110001;
    16'b0010000100000000: out_v[384] = 10'b0111111011;
    16'b0010000110000000: out_v[384] = 10'b0111101111;
    16'b0010010100100100: out_v[384] = 10'b0001011111;
    16'b0010000000000000: out_v[384] = 10'b1000001110;
    16'b0010000101000000: out_v[384] = 10'b1010000101;
    16'b0010000100100000: out_v[384] = 10'b0001011110;
    16'b0010000100101000: out_v[384] = 10'b1100011011;
    16'b0000000100100100: out_v[384] = 10'b1101101100;
    16'b0010100100000110: out_v[384] = 10'b1110110001;
    16'b0010000000000100: out_v[384] = 10'b0110100011;
    16'b0010000100101100: out_v[384] = 10'b0001101110;
    16'b0010100100000000: out_v[384] = 10'b0111001111;
    16'b0000000100100000: out_v[384] = 10'b0110110111;
    16'b0010100100000100: out_v[384] = 10'b1101111110;
    16'b0010000100001100: out_v[384] = 10'b1111001111;
    16'b0010000101100000: out_v[384] = 10'b0110011011;
    16'b0000000000100000: out_v[384] = 10'b0101011011;
    16'b0010110110101100: out_v[384] = 10'b0100011000;
    16'b0010110010001100: out_v[384] = 10'b1011001011;
    16'b0010110110100100: out_v[384] = 10'b0111110000;
    16'b0010010110100100: out_v[384] = 10'b1111110000;
    16'b0000010000100100: out_v[384] = 10'b1111000101;
    16'b0010110110100110: out_v[384] = 10'b0111011011;
    16'b0010110010101100: out_v[384] = 10'b1010100011;
    16'b0000000100001100: out_v[384] = 10'b1101100100;
    16'b1010110111000110: out_v[384] = 10'b1011011010;
    16'b0010000110001100: out_v[384] = 10'b0001001011;
    16'b0010110100000100: out_v[384] = 10'b1001101011;
    16'b0010110100000110: out_v[384] = 10'b1000111111;
    16'b0010010100000000: out_v[384] = 10'b1001011001;
    default: out_v[384] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000110000100000: out_v[385] = 10'b0001010111;
    16'b0000111010100000: out_v[385] = 10'b0000010011;
    16'b0000111010100010: out_v[385] = 10'b0111000111;
    16'b0000100000000000: out_v[385] = 10'b1001010011;
    16'b0100110000100100: out_v[385] = 10'b0011111010;
    16'b1001010000100000: out_v[385] = 10'b0011010101;
    16'b0000010000100010: out_v[385] = 10'b0000111011;
    16'b0100010000100100: out_v[385] = 10'b1000000011;
    16'b0000111000100000: out_v[385] = 10'b1111100011;
    16'b0000111010000000: out_v[385] = 10'b1001111001;
    16'b0000110000100100: out_v[385] = 10'b0001011101;
    16'b1001110000100000: out_v[385] = 10'b1111000110;
    16'b0000110000000000: out_v[385] = 10'b1000010111;
    16'b0000101010000000: out_v[385] = 10'b1000001101;
    16'b0000110010100000: out_v[385] = 10'b1110001001;
    16'b0000111000000000: out_v[385] = 10'b1010011101;
    16'b0001110000100000: out_v[385] = 10'b1000010111;
    16'b1001010000000010: out_v[385] = 10'b1010100110;
    16'b0100111010100000: out_v[385] = 10'b0110101011;
    16'b0000010000100000: out_v[385] = 10'b0010000110;
    16'b0000101000000000: out_v[385] = 10'b0010011001;
    16'b0000011010100000: out_v[385] = 10'b1001110001;
    16'b0001110000000000: out_v[385] = 10'b0010010111;
    16'b1001011010100010: out_v[385] = 10'b0111011010;
    16'b0100111010100100: out_v[385] = 10'b0000100011;
    16'b0001011010100010: out_v[385] = 10'b0101111110;
    16'b1001010000000000: out_v[385] = 10'b0001110110;
    16'b1001110000000000: out_v[385] = 10'b0000110111;
    16'b0000011010100010: out_v[385] = 10'b0011011111;
    16'b0000110010000000: out_v[385] = 10'b1111100110;
    16'b0001011010100000: out_v[385] = 10'b1101010101;
    16'b0000111010100100: out_v[385] = 10'b1100110001;
    16'b0001110010100000: out_v[385] = 10'b1111010100;
    16'b0000110010100100: out_v[385] = 10'b1011011000;
    16'b0100010000000100: out_v[385] = 10'b1100001110;
    16'b0000010000100100: out_v[385] = 10'b0101011100;
    16'b0001111010100000: out_v[385] = 10'b1011010101;
    16'b1001010000100010: out_v[385] = 10'b0011011111;
    16'b0000010010100000: out_v[385] = 10'b0000110101;
    16'b0100010000100000: out_v[385] = 10'b0011001000;
    16'b0000000000100000: out_v[385] = 10'b1110100111;
    16'b0000010000000000: out_v[385] = 10'b1101011100;
    16'b0100000000100000: out_v[385] = 10'b1010001001;
    16'b0000000000000100: out_v[385] = 10'b0011111000;
    16'b0000010000000100: out_v[385] = 10'b0111101000;
    16'b0100001000000100: out_v[385] = 10'b0001010011;
    16'b0000000000000000: out_v[385] = 10'b1011100110;
    16'b0100001010000100: out_v[385] = 10'b1100001011;
    16'b0100000000000100: out_v[385] = 10'b0010110101;
    16'b0000001010000100: out_v[385] = 10'b1001011110;
    16'b0100000000000000: out_v[385] = 10'b1001001100;
    16'b0000001000000000: out_v[385] = 10'b1001101001;
    16'b0000001000000100: out_v[385] = 10'b0100010111;
    16'b0100010000000000: out_v[385] = 10'b1110010000;
    16'b1101010000100100: out_v[385] = 10'b1000100110;
    16'b1101010000000100: out_v[385] = 10'b1111001010;
    16'b0100000010000100: out_v[385] = 10'b1001100011;
    16'b0101010010000100: out_v[385] = 10'b0111100001;
    16'b0100101010000100: out_v[385] = 10'b1011111101;
    16'b1101000010000100: out_v[385] = 10'b0101001101;
    16'b0101000010000100: out_v[385] = 10'b1100001100;
    16'b0101010000000100: out_v[385] = 10'b1011000001;
    16'b1101010010100100: out_v[385] = 10'b0011000111;
    16'b0100000000100100: out_v[385] = 10'b1011100000;
    16'b0100110010000100: out_v[385] = 10'b0101001101;
    16'b1101000000000100: out_v[385] = 10'b0100011011;
    16'b0100010010100100: out_v[385] = 10'b0101001001;
    16'b0100010010000100: out_v[385] = 10'b0100111011;
    16'b1101010010000100: out_v[385] = 10'b0111011001;
    16'b1101001010000100: out_v[385] = 10'b0000011111;
    16'b1001010000000100: out_v[385] = 10'b0100100011;
    16'b0100011010100100: out_v[385] = 10'b0011001100;
    16'b0100011010000100: out_v[385] = 10'b0011011001;
    16'b0100111010000100: out_v[385] = 10'b0010101010;
    16'b0100101010000000: out_v[385] = 10'b1111010100;
    16'b0100110000000100: out_v[385] = 10'b1000110100;
    16'b0100110010100100: out_v[385] = 10'b1001001011;
    16'b1101011010100100: out_v[385] = 10'b1001100011;
    16'b1001010000100100: out_v[385] = 10'b0001001110;
    16'b1101011010000100: out_v[385] = 10'b1010111111;
    16'b0101010000100100: out_v[385] = 10'b0110110100;
    16'b0101000000000100: out_v[385] = 10'b1100000110;
    16'b0101001010000100: out_v[385] = 10'b1110100101;
    16'b0000110010000100: out_v[385] = 10'b1011110111;
    16'b0100010010000000: out_v[385] = 10'b1111010011;
    16'b0000000010000100: out_v[385] = 10'b1010011101;
    16'b0101010000100000: out_v[385] = 10'b0110101000;
    16'b0000101010000100: out_v[385] = 10'b1000111011;
    16'b0101110000100100: out_v[385] = 10'b1001100101;
    16'b0100011000100100: out_v[385] = 10'b1110100000;
    16'b0001110000100100: out_v[385] = 10'b0110111010;
    16'b1101110000100100: out_v[385] = 10'b0111001110;
    16'b1001110000100100: out_v[385] = 10'b0100001011;
    16'b0000011010000100: out_v[385] = 10'b1011011110;
    16'b0000100010000100: out_v[385] = 10'b1011110100;
    16'b0000010010000100: out_v[385] = 10'b1111111011;
    16'b0001110010000100: out_v[385] = 10'b1111100010;
    16'b0000110000000100: out_v[385] = 10'b1110100011;
    16'b0001110010100100: out_v[385] = 10'b0110011101;
    16'b0000111010000100: out_v[385] = 10'b0001001010;
    16'b1101110010100100: out_v[385] = 10'b1100001110;
    16'b1101010000100000: out_v[385] = 10'b0111001010;
    16'b0000010010100100: out_v[385] = 10'b0100001101;
    16'b0100100000000100: out_v[385] = 10'b0011111000;
    16'b0100101000000100: out_v[385] = 10'b0000110000;
    16'b0101100000000100: out_v[385] = 10'b1100001011;
    16'b0100001000100100: out_v[385] = 10'b0000011011;
    16'b0100101000000000: out_v[385] = 10'b0100011011;
    16'b1101100000000100: out_v[385] = 10'b0001111011;
    16'b0100100000000000: out_v[385] = 10'b0101011110;
    16'b0100100000100100: out_v[385] = 10'b1010100111;
    16'b0100000010000000: out_v[385] = 10'b1010111000;
    16'b0100011000100000: out_v[385] = 10'b1010100001;
    16'b0100011000000100: out_v[385] = 10'b1110000011;
    16'b0100001010100000: out_v[385] = 10'b1010101100;
    16'b0000011000100000: out_v[385] = 10'b0001110010;
    16'b0100001000100000: out_v[385] = 10'b1001010111;
    16'b0000001000100000: out_v[385] = 10'b0001111110;
    16'b0100011010100000: out_v[385] = 10'b0110010101;
    16'b1001100000000100: out_v[385] = 10'b1011001010;
    16'b1001110000000100: out_v[385] = 10'b0010011010;
    16'b0100010010100000: out_v[385] = 10'b0010101110;
    16'b0001110000000100: out_v[385] = 10'b0100111010;
    16'b0100011000000000: out_v[385] = 10'b0111010001;
    16'b0000100000000100: out_v[385] = 10'b1011001010;
    16'b0000001010000000: out_v[385] = 10'b0001001100;
    16'b0101011000100000: out_v[385] = 10'b0010111001;
    16'b0000000010000000: out_v[385] = 10'b1010110110;
    16'b0100001010000000: out_v[385] = 10'b1111001110;
    16'b0000111000100100: out_v[385] = 10'b1010100000;
    16'b0000011010100100: out_v[385] = 10'b0111001110;
    16'b0100001000000000: out_v[385] = 10'b1101101000;
    16'b0001100000000100: out_v[385] = 10'b1010111010;
    16'b0100000000000110: out_v[385] = 10'b0101100010;
    16'b0100110000100000: out_v[385] = 10'b1101000110;
    16'b0100100000000110: out_v[385] = 10'b0000011100;
    16'b0100111000100100: out_v[385] = 10'b1010000011;
    16'b0000100000100100: out_v[385] = 10'b1110011010;
    16'b0100100000100000: out_v[385] = 10'b1111000111;
    16'b0000100000100000: out_v[385] = 10'b0101010101;
    16'b0000000000100100: out_v[385] = 10'b1100001101;
    16'b0100101000100100: out_v[385] = 10'b0011001111;
    16'b0000011000000100: out_v[385] = 10'b0011011011;
    16'b0000011000100100: out_v[385] = 10'b1111111100;
    default: out_v[385] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0101000000001000: out_v[386] = 10'b1100101101;
    16'b0000000100001010: out_v[386] = 10'b0101010001;
    16'b0001000100001010: out_v[386] = 10'b0100010011;
    16'b0001000000000000: out_v[386] = 10'b1011011010;
    16'b0100000000001000: out_v[386] = 10'b1011000101;
    16'b0001000000001000: out_v[386] = 10'b1110110000;
    16'b0000000000001000: out_v[386] = 10'b0001011110;
    16'b0000000000000000: out_v[386] = 10'b0111001101;
    16'b1000000100001010: out_v[386] = 10'b0010000011;
    16'b0001010000001000: out_v[386] = 10'b0000110011;
    16'b0101010000001000: out_v[386] = 10'b1000111001;
    16'b1000000000001000: out_v[386] = 10'b0100110001;
    16'b0100000100001010: out_v[386] = 10'b0110111001;
    16'b1001000100001010: out_v[386] = 10'b1010010011;
    16'b0001010000000000: out_v[386] = 10'b1101001000;
    16'b0101000100001010: out_v[386] = 10'b0000100110;
    16'b1001000000001000: out_v[386] = 10'b0000110010;
    16'b1001010000001000: out_v[386] = 10'b0001101001;
    16'b0001010000001100: out_v[386] = 10'b1111100001;
    16'b0100000000000000: out_v[386] = 10'b0011111010;
    16'b0000000100000010: out_v[386] = 10'b1100101100;
    16'b0001010100001010: out_v[386] = 10'b0010100010;
    16'b0101000000000000: out_v[386] = 10'b0011010100;
    16'b0000010000001000: out_v[386] = 10'b0011100100;
    16'b0100000100000010: out_v[386] = 10'b1010001011;
    16'b0001000000001100: out_v[386] = 10'b0001011110;
    16'b0000010000000000: out_v[386] = 10'b1111000100;
    16'b0101000100000010: out_v[386] = 10'b1110010011;
    16'b0000010100001010: out_v[386] = 10'b1111010111;
    16'b0100010000001000: out_v[386] = 10'b0010010011;
    16'b0101010000001100: out_v[386] = 10'b0001110101;
    16'b0100000000001100: out_v[386] = 10'b1010001110;
    16'b0100010100001110: out_v[386] = 10'b0010110111;
    16'b0101010100001010: out_v[386] = 10'b1000011010;
    16'b0100010000000000: out_v[386] = 10'b1001001011;
    16'b0100000100001110: out_v[386] = 10'b1011110010;
    16'b0100010000001100: out_v[386] = 10'b1011011110;
    16'b0100010100001010: out_v[386] = 10'b1010011000;
    16'b0101000000001100: out_v[386] = 10'b0010010110;
    16'b0101010100001110: out_v[386] = 10'b1101110110;
    16'b0100010100000010: out_v[386] = 10'b0111110110;
    16'b0000000000001100: out_v[386] = 10'b0000101110;
    16'b0100000010001000: out_v[386] = 10'b0010001010;
    16'b0101010100000010: out_v[386] = 10'b1111101010;
    16'b0101010000000000: out_v[386] = 10'b0100111000;
    16'b0001010100000010: out_v[386] = 10'b1000011110;
    16'b0001000100000010: out_v[386] = 10'b1001000110;
    16'b1100000000000000: out_v[386] = 10'b1011000111;
    16'b0100010000000100: out_v[386] = 10'b1000011110;
    16'b1000000100000010: out_v[386] = 10'b1011100111;
    16'b1000000000000000: out_v[386] = 10'b0000101000;
    16'b0000001000001000: out_v[386] = 10'b0100100001;
    16'b0100001000001000: out_v[386] = 10'b0011100010;
    16'b0000001000000000: out_v[386] = 10'b0101000100;
    16'b0100001000000000: out_v[386] = 10'b0101001110;
    16'b1100000100001010: out_v[386] = 10'b0101010000;
    16'b1100000000001000: out_v[386] = 10'b1100010001;
    16'b1101000000001000: out_v[386] = 10'b0110001110;
    16'b1101000100001010: out_v[386] = 10'b0101010000;
    16'b1101010000001000: out_v[386] = 10'b0101000010;
    default: out_v[386] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b1000100001000000: out_v[387] = 10'b1001011101;
    16'b1000100101110101: out_v[387] = 10'b0010110001;
    16'b1000100101000000: out_v[387] = 10'b0111010001;
    16'b0000000100100000: out_v[387] = 10'b1011101000;
    16'b1000100100100000: out_v[387] = 10'b0100100101;
    16'b0000000100110101: out_v[387] = 10'b0011011111;
    16'b1000100100110001: out_v[387] = 10'b0100110111;
    16'b0000000100000000: out_v[387] = 10'b1001011011;
    16'b0000100101110001: out_v[387] = 10'b1110010110;
    16'b1000100101110001: out_v[387] = 10'b0110001101;
    16'b1000100001000001: out_v[387] = 10'b0001101011;
    16'b1000100101100001: out_v[387] = 10'b0001011011;
    16'b1000100101010001: out_v[387] = 10'b1100111010;
    16'b0000100101010101: out_v[387] = 10'b1101011011;
    16'b0000000100110000: out_v[387] = 10'b1001110010;
    16'b1000100101100000: out_v[387] = 10'b0101000000;
    16'b0000000100110001: out_v[387] = 10'b0101000011;
    16'b1000000100100000: out_v[387] = 10'b1001001110;
    16'b0000100101100000: out_v[387] = 10'b1111000100;
    16'b0000100101110101: out_v[387] = 10'b1010110110;
    16'b1000100101010101: out_v[387] = 10'b0100010001;
    16'b1000100101000001: out_v[387] = 10'b1101000011;
    16'b0000000000110101: out_v[387] = 10'b0101101011;
    16'b1000100101000101: out_v[387] = 10'b1000000111;
    16'b1000100101110000: out_v[387] = 10'b1111000011;
    16'b0000000101110001: out_v[387] = 10'b1011011110;
    16'b0000000101110101: out_v[387] = 10'b1111011100;
    16'b1000100101000100: out_v[387] = 10'b1101110111;
    16'b0000000100100001: out_v[387] = 10'b1111011011;
    16'b1000000100110001: out_v[387] = 10'b1111000101;
    16'b1000100001100000: out_v[387] = 10'b0001001010;
    16'b1000100101100101: out_v[387] = 10'b1110000111;
    16'b0000000001110101: out_v[387] = 10'b1001001111;
    16'b1000100101100100: out_v[387] = 10'b0111100011;
    16'b0000000000000000: out_v[387] = 10'b0101000111;
    16'b1000000000000000: out_v[387] = 10'b1110001000;
    16'b0000000000000001: out_v[387] = 10'b1101000011;
    16'b0000000000000100: out_v[387] = 10'b0000011111;
    16'b1000000000000101: out_v[387] = 10'b0101010110;
    16'b1000000000000001: out_v[387] = 10'b1011000101;
    16'b1000000100000101: out_v[387] = 10'b0110010100;
    16'b0000000000000101: out_v[387] = 10'b0000101111;
    16'b0000000001000000: out_v[387] = 10'b1101000001;
    16'b0000000000000010: out_v[387] = 10'b0000001111;
    16'b1000000100000001: out_v[387] = 10'b0010111101;
    16'b1000000100000000: out_v[387] = 10'b1011101100;
    16'b1000100100000000: out_v[387] = 10'b0111100100;
    16'b0000100101000000: out_v[387] = 10'b1000110100;
    16'b1000000100000100: out_v[387] = 10'b0100100100;
    16'b1000100000000000: out_v[387] = 10'b1001001010;
    16'b0000100100000000: out_v[387] = 10'b0110000110;
    16'b1000100100000100: out_v[387] = 10'b1101011000;
    16'b1000100100000010: out_v[387] = 10'b0111000111;
    16'b1000100101000010: out_v[387] = 10'b0110000110;
    16'b1000000100000110: out_v[387] = 10'b1101110011;
    16'b1000000100000010: out_v[387] = 10'b1001101011;
    16'b1000100100000101: out_v[387] = 10'b1001110111;
    16'b1000000100010101: out_v[387] = 10'b0010010111;
    16'b1000000000000010: out_v[387] = 10'b1000110111;
    16'b1000100000000010: out_v[387] = 10'b1110111010;
    16'b1000100100000001: out_v[387] = 10'b0100100111;
    16'b1000100100010101: out_v[387] = 10'b1111000110;
    16'b1000000000000100: out_v[387] = 10'b0100010011;
    16'b1000100100010001: out_v[387] = 10'b0111000111;
    16'b1000000100000111: out_v[387] = 10'b1000111011;
    16'b0000000001000100: out_v[387] = 10'b1011110100;
    16'b0000000101000100: out_v[387] = 10'b0011110100;
    16'b0000000001010101: out_v[387] = 10'b1101001001;
    16'b0000100001000100: out_v[387] = 10'b0010100011;
    16'b0000000000010101: out_v[387] = 10'b0000111011;
    16'b0000000001100000: out_v[387] = 10'b0100100100;
    16'b0000100001000010: out_v[387] = 10'b1000011011;
    16'b0000000001000010: out_v[387] = 10'b0101110011;
    16'b0000100001000000: out_v[387] = 10'b0010101000;
    16'b0000000100000101: out_v[387] = 10'b1011100011;
    16'b0000100001100100: out_v[387] = 10'b0011001110;
    16'b0000100001000101: out_v[387] = 10'b1001001110;
    16'b0000000101000000: out_v[387] = 10'b1011001111;
    16'b0000000001000101: out_v[387] = 10'b1101010110;
    16'b0000100000000000: out_v[387] = 10'b1110000000;
    16'b0000000100000001: out_v[387] = 10'b1010111000;
    16'b0000100001010101: out_v[387] = 10'b1011111100;
    16'b0000100001100000: out_v[387] = 10'b0010111010;
    16'b0000000001100100: out_v[387] = 10'b0100011111;
    16'b1000000101000000: out_v[387] = 10'b0010101100;
    16'b0000000100000100: out_v[387] = 10'b0011101100;
    16'b1000100000000001: out_v[387] = 10'b1100011010;
    16'b0000100001010001: out_v[387] = 10'b0011011011;
    16'b0000100001000001: out_v[387] = 10'b0110110001;
    16'b1000100000010001: out_v[387] = 10'b1101100000;
    16'b0000000001000001: out_v[387] = 10'b0111110111;
    16'b1000100001010001: out_v[387] = 10'b0111001010;
    16'b1000100000100000: out_v[387] = 10'b1011000001;
    16'b0000100000000001: out_v[387] = 10'b1111111110;
    16'b1000100001100001: out_v[387] = 10'b0000111101;
    16'b0000100001010000: out_v[387] = 10'b0011110000;
    16'b0000100001100001: out_v[387] = 10'b1101110100;
    16'b1000100001010000: out_v[387] = 10'b0010111010;
    16'b0000000101010001: out_v[387] = 10'b1011111110;
    16'b0000000001010000: out_v[387] = 10'b0001100111;
    16'b0000000101000001: out_v[387] = 10'b0000100110;
    16'b0000100101000001: out_v[387] = 10'b0100101011;
    16'b0000100101010001: out_v[387] = 10'b1010111010;
    16'b0000100101010000: out_v[387] = 10'b1000001101;
    16'b0000100101000101: out_v[387] = 10'b1010101111;
    16'b1000000101000001: out_v[387] = 10'b1010101110;
    16'b1000100001000101: out_v[387] = 10'b1010111000;
    16'b0000000101010000: out_v[387] = 10'b0001110110;
    16'b0000000001010001: out_v[387] = 10'b1111010010;
    16'b0000000101000101: out_v[387] = 10'b1011101011;
    16'b1000000001000000: out_v[387] = 10'b0110100110;
    16'b0000000000010001: out_v[387] = 10'b0111001110;
    16'b0000001000000001: out_v[387] = 10'b0111110010;
    16'b0000001000010001: out_v[387] = 10'b0101011101;
    16'b0100000000000000: out_v[387] = 10'b0110010010;
    16'b0000000000100000: out_v[387] = 10'b0110000111;
    16'b0000000000010000: out_v[387] = 10'b1110100110;
    16'b0100000000010000: out_v[387] = 10'b0011111101;
    16'b0000001000010000: out_v[387] = 10'b0111111011;
    16'b0000001000000000: out_v[387] = 10'b0101110101;
    16'b0000001001010001: out_v[387] = 10'b0111000011;
    16'b1000000101010101: out_v[387] = 10'b0011111010;
    16'b1000000001000001: out_v[387] = 10'b1000110100;
    16'b1000000000010000: out_v[387] = 10'b1100010101;
    16'b1000000000010001: out_v[387] = 10'b0110011011;
    16'b1000000000010101: out_v[387] = 10'b1100010011;
    16'b1000000001010001: out_v[387] = 10'b0000001110;
    16'b1000100001000010: out_v[387] = 10'b0111010110;
    16'b1000000001010000: out_v[387] = 10'b0100011011;
    default: out_v[387] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000001000000000: out_v[388] = 10'b1011111011;
    16'b0000001000011000: out_v[388] = 10'b1000010001;
    16'b1000001000011000: out_v[388] = 10'b0010000011;
    16'b1000011000011000: out_v[388] = 10'b0001000001;
    16'b0000000000001000: out_v[388] = 10'b0000101110;
    16'b0000011000011000: out_v[388] = 10'b0001010000;
    16'b0000000000011000: out_v[388] = 10'b0101101011;
    16'b1000000000001000: out_v[388] = 10'b1100110101;
    16'b0000010000011000: out_v[388] = 10'b1010011110;
    16'b1000010000011000: out_v[388] = 10'b0101100011;
    16'b0000001000010000: out_v[388] = 10'b1010011011;
    16'b1000001000010000: out_v[388] = 10'b1111010110;
    16'b1000001000001000: out_v[388] = 10'b1010100110;
    16'b0000000000010000: out_v[388] = 10'b0100100011;
    16'b1000000000011000: out_v[388] = 10'b0111000101;
    16'b0000001000001000: out_v[388] = 10'b1001000101;
    16'b0000000000000000: out_v[388] = 10'b0110001011;
    16'b1000000000010000: out_v[388] = 10'b1001001011;
    16'b0000010000001000: out_v[388] = 10'b1100000110;
    16'b1000000000000000: out_v[388] = 10'b0101001011;
    16'b1000010000001000: out_v[388] = 10'b0110011010;
    16'b0000010000000000: out_v[388] = 10'b1100010100;
    16'b1000010000000000: out_v[388] = 10'b0101100100;
    16'b0001000000001000: out_v[388] = 10'b1011000100;
    16'b0001010000001000: out_v[388] = 10'b1110100100;
    16'b0000010000010000: out_v[388] = 10'b1100010100;
    16'b1001000000001000: out_v[388] = 10'b1100001100;
    16'b1000011000001000: out_v[388] = 10'b1010111011;
    16'b0000011000010000: out_v[388] = 10'b1100100000;
    16'b1000010000010000: out_v[388] = 10'b1010001110;
    16'b0000011000001000: out_v[388] = 10'b1111101100;
    16'b1001010000001000: out_v[388] = 10'b1101010011;
    16'b0000011000000000: out_v[388] = 10'b0111111010;
    16'b1000011000010000: out_v[388] = 10'b0111010010;
    16'b0001011000001000: out_v[388] = 10'b0110001100;
    16'b0001010000011000: out_v[388] = 10'b0110011011;
    16'b0001001000001000: out_v[388] = 10'b1111111010;
    16'b1000011000000000: out_v[388] = 10'b0101111100;
    16'b0001010000000000: out_v[388] = 10'b0111011010;
    16'b0001011000000000: out_v[388] = 10'b1011001000;
    16'b1001011000001000: out_v[388] = 10'b0110110000;
    16'b0001000000000000: out_v[388] = 10'b1011111100;
    16'b0001011000011000: out_v[388] = 10'b1101110111;
    16'b0001001000000000: out_v[388] = 10'b1000110110;
    16'b0001011000010000: out_v[388] = 10'b0000111011;
    16'b0010011000000000: out_v[388] = 10'b0011101111;
    16'b0000010001011000: out_v[388] = 10'b0010111100;
    16'b0000010001010000: out_v[388] = 10'b1100010010;
    16'b0001010000010000: out_v[388] = 10'b1101101011;
    16'b0000000001001000: out_v[388] = 10'b1000111011;
    16'b0000000001000000: out_v[388] = 10'b1100011000;
    16'b0000000001010000: out_v[388] = 10'b0000100110;
    16'b0000000001011000: out_v[388] = 10'b1000101010;
    16'b0000010001001000: out_v[388] = 10'b0100001101;
    16'b1000001000000000: out_v[388] = 10'b1001100100;
    16'b0001000000011000: out_v[388] = 10'b1011011001;
    16'b0001001000011000: out_v[388] = 10'b1011010011;
    16'b0010011000001000: out_v[388] = 10'b0111001000;
    16'b0010010000001000: out_v[388] = 10'b0010101010;
    16'b0010010000000000: out_v[388] = 10'b0110011011;
    16'b0010001000001000: out_v[388] = 10'b1111111000;
    16'b0010001000000000: out_v[388] = 10'b1011010011;
    16'b0000010000000010: out_v[388] = 10'b1011110010;
    16'b0000010001000000: out_v[388] = 10'b1101001011;
    default: out_v[388] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000001001000000: out_v[389] = 10'b0000000111;
    16'b0000000001000000: out_v[389] = 10'b0010110101;
    16'b1000001100000000: out_v[389] = 10'b1110001111;
    16'b1000001000000000: out_v[389] = 10'b1110011011;
    16'b0000001001000100: out_v[389] = 10'b0000111011;
    16'b0000001000000000: out_v[389] = 10'b0000111100;
    16'b1000000000000000: out_v[389] = 10'b0000010001;
    16'b1000001001000000: out_v[389] = 10'b0100000111;
    16'b0000000001000001: out_v[389] = 10'b1010110101;
    16'b1000001101000000: out_v[389] = 10'b0110001111;
    16'b0000000001000100: out_v[389] = 10'b0111011100;
    16'b1000000001000000: out_v[389] = 10'b0110000000;
    16'b0000001001000101: out_v[389] = 10'b0011100011;
    16'b1000000100000000: out_v[389] = 10'b1111011110;
    16'b0000001001000001: out_v[389] = 10'b1001010111;
    16'b0000000000000000: out_v[389] = 10'b0001101000;
    16'b1000001010000000: out_v[389] = 10'b1100100011;
    16'b1000001011000000: out_v[389] = 10'b0000110001;
    16'b1000000101000000: out_v[389] = 10'b1111011011;
    16'b1000001001000001: out_v[389] = 10'b1010110011;
    16'b0000001001001001: out_v[389] = 10'b1111010110;
    16'b0001001000001101: out_v[389] = 10'b0010001010;
    16'b0001000000001101: out_v[389] = 10'b1000011011;
    16'b0001000000001001: out_v[389] = 10'b0110011100;
    16'b0000000000001001: out_v[389] = 10'b0111001000;
    16'b0000000000000001: out_v[389] = 10'b1000100111;
    16'b0000001000001001: out_v[389] = 10'b0001001100;
    16'b0001000000000101: out_v[389] = 10'b0101111001;
    16'b0001000000001100: out_v[389] = 10'b0010010101;
    16'b0001001000001001: out_v[389] = 10'b1001101111;
    16'b0001000000001000: out_v[389] = 10'b1111001001;
    16'b0001000000000001: out_v[389] = 10'b1101110011;
    16'b0000000000001000: out_v[389] = 10'b1110001011;
    16'b0001001000001100: out_v[389] = 10'b0110010011;
    16'b0001001001000101: out_v[389] = 10'b0011000101;
    16'b0001000000000100: out_v[389] = 10'b0011001110;
    16'b0001001000000100: out_v[389] = 10'b0011000100;
    16'b0000001010000100: out_v[389] = 10'b0111100010;
    16'b0001000001000101: out_v[389] = 10'b0010111100;
    16'b0000000010001001: out_v[389] = 10'b1001011101;
    16'b0001000001000100: out_v[389] = 10'b1100010100;
    16'b0001001001001101: out_v[389] = 10'b0010101110;
    16'b0000001000000100: out_v[389] = 10'b1011000100;
    16'b0001001010000100: out_v[389] = 10'b1000010011;
    16'b0000000000000100: out_v[389] = 10'b0110010100;
    16'b0001001001000100: out_v[389] = 10'b1111001000;
    16'b0001001001001100: out_v[389] = 10'b1010110001;
    16'b0001000010000100: out_v[389] = 10'b1000011000;
    16'b0000000001001001: out_v[389] = 10'b1001101100;
    16'b0000001010000000: out_v[389] = 10'b0010010110;
    16'b0001000001001101: out_v[389] = 10'b0010001011;
    16'b0001001010001100: out_v[389] = 10'b1111110001;
    16'b0001001000000101: out_v[389] = 10'b1100110001;
    16'b0001000010001100: out_v[389] = 10'b0010100101;
    16'b0001001010001101: out_v[389] = 10'b0100001011;
    16'b0000001010001001: out_v[389] = 10'b1011001011;
    16'b0001000011000101: out_v[389] = 10'b0111101011;
    16'b0000001000001101: out_v[389] = 10'b0010101010;
    16'b0000000010001101: out_v[389] = 10'b1111011001;
    16'b0000000000001101: out_v[389] = 10'b1101000000;
    16'b0000000001001101: out_v[389] = 10'b1101100010;
    16'b0001000010000101: out_v[389] = 10'b0100001011;
    16'b0001000010001101: out_v[389] = 10'b1111110011;
    16'b0001000011001101: out_v[389] = 10'b0000011011;
    16'b0000001001001101: out_v[389] = 10'b0111110100;
    16'b0000000000001100: out_v[389] = 10'b1010101001;
    16'b0000000000000101: out_v[389] = 10'b1001001001;
    16'b0000001000001000: out_v[389] = 10'b0100111001;
    16'b0000000011001001: out_v[389] = 10'b1100101010;
    16'b0001000001001100: out_v[389] = 10'b0100110011;
    16'b0001000101000101: out_v[389] = 10'b0011110001;
    16'b0001000101000100: out_v[389] = 10'b1100110011;
    16'b1001000001001101: out_v[389] = 10'b0000010100;
    16'b1001000001000100: out_v[389] = 10'b1100011010;
    16'b0001000011000100: out_v[389] = 10'b1010101010;
    16'b1001000001001100: out_v[389] = 10'b1010110010;
    16'b0000000001000101: out_v[389] = 10'b0010110101;
    16'b0001000001010100: out_v[389] = 10'b1111001011;
    16'b1001000001000101: out_v[389] = 10'b0111010110;
    16'b0000001100000000: out_v[389] = 10'b0100011111;
    16'b0001001101000101: out_v[389] = 10'b1011110000;
    16'b0001001100000101: out_v[389] = 10'b1011010110;
    16'b0001001100001101: out_v[389] = 10'b1101110111;
    16'b0001000100000101: out_v[389] = 10'b1011011111;
    16'b0000001000000001: out_v[389] = 10'b0010100110;
    16'b0000000101000000: out_v[389] = 10'b1001100010;
    16'b0000001101000000: out_v[389] = 10'b1011011011;
    16'b0001001101000100: out_v[389] = 10'b0100111011;
    16'b0000001000000101: out_v[389] = 10'b0000111011;
    16'b0000000100000000: out_v[389] = 10'b0000110010;
    16'b0001001001100100: out_v[389] = 10'b1110010000;
    16'b0001001001100101: out_v[389] = 10'b1110010111;
    16'b1001001001000100: out_v[389] = 10'b1001011100;
    16'b1001001001100100: out_v[389] = 10'b0011110101;
    16'b1001000000000100: out_v[389] = 10'b1001101100;
    16'b0001000001100100: out_v[389] = 10'b1010101111;
    16'b0001000000100100: out_v[389] = 10'b0111011011;
    16'b1001001001000101: out_v[389] = 10'b1001110010;
    16'b1000000001001001: out_v[389] = 10'b0011101110;
    16'b0001000001100101: out_v[389] = 10'b0110001011;
    16'b0001000000100101: out_v[389] = 10'b1110110011;
    16'b1001001000000100: out_v[389] = 10'b0111100110;
    16'b1000001001001001: out_v[389] = 10'b1011111010;
    16'b1001001001001101: out_v[389] = 10'b1010110110;
    16'b0000000001100100: out_v[389] = 10'b1101101110;
    16'b0000000010000000: out_v[389] = 10'b0010110100;
    16'b0000000010000100: out_v[389] = 10'b1000001111;
    16'b0001000100000100: out_v[389] = 10'b1110100111;
    16'b0001001000000001: out_v[389] = 10'b1010100011;
    16'b0001000100001101: out_v[389] = 10'b0111010101;
    16'b0001000101001101: out_v[389] = 10'b0111001010;
    16'b0001001100000100: out_v[389] = 10'b1111001000;
    16'b0001001101001101: out_v[389] = 10'b1001101010;
    default: out_v[389] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0001010000010100: out_v[390] = 10'b0000110011;
    16'b1000011000010000: out_v[390] = 10'b1110100001;
    16'b1101011000010100: out_v[390] = 10'b0000001001;
    16'b1100010000010100: out_v[390] = 10'b1111101011;
    16'b1000010000010100: out_v[390] = 10'b1101011000;
    16'b0101010001000100: out_v[390] = 10'b1100011111;
    16'b1101010000000100: out_v[390] = 10'b0111000010;
    16'b0100010000000000: out_v[390] = 10'b0100110001;
    16'b0000000000000100: out_v[390] = 10'b0001100011;
    16'b1001010000000100: out_v[390] = 10'b1100010100;
    16'b1101010000010100: out_v[390] = 10'b0001100001;
    16'b1001011010010100: out_v[390] = 10'b0101001001;
    16'b1000010000010000: out_v[390] = 10'b1111100111;
    16'b0000010000010100: out_v[390] = 10'b1100110001;
    16'b0000010000010000: out_v[390] = 10'b1111110011;
    16'b1000010000000100: out_v[390] = 10'b1000111011;
    16'b1001010000010100: out_v[390] = 10'b1100010100;
    16'b0101010000010100: out_v[390] = 10'b0111000001;
    16'b0100010000010100: out_v[390] = 10'b0011011011;
    16'b1000011000010100: out_v[390] = 10'b1001011110;
    16'b0101010000000100: out_v[390] = 10'b0111011111;
    16'b0001000000010100: out_v[390] = 10'b0010001101;
    16'b0100010000000100: out_v[390] = 10'b1111011101;
    16'b0100100001000100: out_v[390] = 10'b1001100111;
    16'b1001011000010100: out_v[390] = 10'b0110001011;
    16'b0100000000000000: out_v[390] = 10'b0100110110;
    16'b0000011000010000: out_v[390] = 10'b0100011110;
    16'b1000011000000100: out_v[390] = 10'b1101010111;
    16'b1001011000000100: out_v[390] = 10'b1100100001;
    16'b0000000000010100: out_v[390] = 10'b0011100111;
    16'b1100010000010000: out_v[390] = 10'b0010011000;
    16'b0100100001000000: out_v[390] = 10'b1011010011;
    16'b1000011010010100: out_v[390] = 10'b0011110101;
    16'b0101110001000100: out_v[390] = 10'b0000010111;
    16'b0100010000010000: out_v[390] = 10'b0011011011;
    16'b0000010000000100: out_v[390] = 10'b1101101011;
    16'b0100000000010000: out_v[390] = 10'b0011011011;
    16'b1001011010000100: out_v[390] = 10'b0011011001;
    16'b1101000000010100: out_v[390] = 10'b1101011001;
    16'b0100000000010100: out_v[390] = 10'b1101101101;
    16'b0100010001000100: out_v[390] = 10'b0010001111;
    16'b1100011000010100: out_v[390] = 10'b1110111100;
    16'b1101011010010100: out_v[390] = 10'b0001101011;
    16'b0000000000010000: out_v[390] = 10'b1011100111;
    16'b0100000000000100: out_v[390] = 10'b1101001110;
    16'b0001001010000100: out_v[390] = 10'b1000010010;
    16'b0000001010000000: out_v[390] = 10'b1100100100;
    16'b0000011010000000: out_v[390] = 10'b1100001010;
    16'b0001000000000000: out_v[390] = 10'b1001011100;
    16'b1000011010000000: out_v[390] = 10'b0000111101;
    16'b0001001010000000: out_v[390] = 10'b1100110010;
    16'b0001000010000100: out_v[390] = 10'b1000000111;
    16'b0000000000000000: out_v[390] = 10'b0010110011;
    16'b1001001010000100: out_v[390] = 10'b1001100011;
    16'b0001000000000100: out_v[390] = 10'b0111001011;
    16'b0000001000000000: out_v[390] = 10'b1010011000;
    16'b1001001010000000: out_v[390] = 10'b0100110010;
    16'b0001000010000000: out_v[390] = 10'b0111001001;
    16'b1000001010000000: out_v[390] = 10'b0101100001;
    16'b1000011000000000: out_v[390] = 10'b0010100110;
    16'b1001011010000000: out_v[390] = 10'b0011010001;
    16'b0000000010000000: out_v[390] = 10'b1011010100;
    16'b0001010000000100: out_v[390] = 10'b1001010110;
    16'b1001111010000100: out_v[390] = 10'b0000100101;
    16'b1001000000000100: out_v[390] = 10'b1010110111;
    16'b1001000010000100: out_v[390] = 10'b1100001100;
    16'b0001111010000100: out_v[390] = 10'b1001111110;
    16'b1001110000000100: out_v[390] = 10'b1100000011;
    16'b1001100000000100: out_v[390] = 10'b0001011100;
    16'b0001011010000100: out_v[390] = 10'b1110000110;
    16'b1001000000010100: out_v[390] = 10'b1100000000;
    16'b1001000001010100: out_v[390] = 10'b1101111101;
    16'b1000000000000000: out_v[390] = 10'b0010111001;
    16'b0001010010000100: out_v[390] = 10'b1001010101;
    16'b1001011011000100: out_v[390] = 10'b0110010101;
    16'b0001110000000100: out_v[390] = 10'b1111000100;
    16'b1000000000000100: out_v[390] = 10'b0010101100;
    16'b1001010001000100: out_v[390] = 10'b1001110011;
    16'b1001110010000100: out_v[390] = 10'b0111110011;
    16'b1000010000000000: out_v[390] = 10'b0111011000;
    16'b1001000000000000: out_v[390] = 10'b1000110100;
    16'b1001010010000100: out_v[390] = 10'b0110110001;
    16'b1001111011000100: out_v[390] = 10'b1011000101;
    16'b0001110010000100: out_v[390] = 10'b1011111110;
    16'b1001110000010100: out_v[390] = 10'b0000001110;
    16'b1001000001000100: out_v[390] = 10'b0100011010;
    16'b0000011010010000: out_v[390] = 10'b0110110001;
    16'b1000011010000100: out_v[390] = 10'b1011111000;
    16'b0001011010010100: out_v[390] = 10'b1000111010;
    16'b1000011010010000: out_v[390] = 10'b1000011100;
    16'b0000001010010000: out_v[390] = 10'b0100001111;
    16'b0000011010000100: out_v[390] = 10'b0111011011;
    16'b0000101010010100: out_v[390] = 10'b0011111011;
    16'b0000001010000100: out_v[390] = 10'b0111000001;
    16'b1000010010000100: out_v[390] = 10'b1100001001;
    16'b0000001010010100: out_v[390] = 10'b0101011110;
    16'b0001001010010100: out_v[390] = 10'b1000011010;
    16'b1000010010000000: out_v[390] = 10'b0000111101;
    16'b0000011010010100: out_v[390] = 10'b1001000000;
    16'b0000101010010000: out_v[390] = 10'b1111011111;
    16'b0000011000000000: out_v[390] = 10'b1000011110;
    16'b1001010000000000: out_v[390] = 10'b1011101010;
    16'b1100000000000000: out_v[390] = 10'b1010110011;
    16'b1100010000100000: out_v[390] = 10'b1111000011;
    16'b0101000000000100: out_v[390] = 10'b1111001010;
    16'b1100010000000000: out_v[390] = 10'b0001011110;
    16'b1100010010010000: out_v[390] = 10'b1001010111;
    16'b1100011010010000: out_v[390] = 10'b1110001110;
    16'b1000000010000000: out_v[390] = 10'b1101001011;
    16'b1100010010000000: out_v[390] = 10'b0000111011;
    16'b1000000000010000: out_v[390] = 10'b0010011000;
    16'b1000010010100000: out_v[390] = 10'b0101110111;
    16'b0001001000000100: out_v[390] = 10'b0110010011;
    16'b1000010000100000: out_v[390] = 10'b0111010111;
    16'b0101000000010100: out_v[390] = 10'b1010010000;
    16'b1100011010000000: out_v[390] = 10'b0001100110;
    16'b1000011010100000: out_v[390] = 10'b1101000100;
    16'b1101010000010000: out_v[390] = 10'b1000011101;
    16'b1101000000010000: out_v[390] = 10'b0100010011;
    16'b1100000000010000: out_v[390] = 10'b1100001110;
    16'b1000001000000000: out_v[390] = 10'b1001001111;
    16'b1000001010000100: out_v[390] = 10'b1101000000;
    16'b1001001000000100: out_v[390] = 10'b0111001101;
    16'b0000010010000000: out_v[390] = 10'b1011100101;
    16'b0000010000000000: out_v[390] = 10'b0100111100;
    16'b0001011000010100: out_v[390] = 10'b1101101000;
    16'b0001010000010000: out_v[390] = 10'b0001011111;
    16'b1001010010010100: out_v[390] = 10'b1000100111;
    16'b1001010000010000: out_v[390] = 10'b0001101110;
    16'b1101010001000100: out_v[390] = 10'b0111011010;
    16'b0001011010000000: out_v[390] = 10'b1111000101;
    16'b0001011000000100: out_v[390] = 10'b0010100100;
    16'b1001001000010100: out_v[390] = 10'b1001100010;
    16'b1001011000010110: out_v[390] = 10'b0111101010;
    16'b0001010000000000: out_v[390] = 10'b0100111100;
    16'b0001011010010000: out_v[390] = 10'b0001011011;
    16'b1001011010000110: out_v[390] = 10'b0001111111;
    16'b1101010001010100: out_v[390] = 10'b1110000101;
    16'b0001010010010100: out_v[390] = 10'b0110101010;
    16'b1000011000100000: out_v[390] = 10'b1001100010;
    16'b1000010000110000: out_v[390] = 10'b0111110100;
    16'b1000011000110000: out_v[390] = 10'b0010001111;
    16'b1000010000100001: out_v[390] = 10'b1110011010;
    16'b1100010000110000: out_v[390] = 10'b0110011110;
    16'b1100011000000000: out_v[390] = 10'b0110001101;
    16'b1001010000100000: out_v[390] = 10'b1001101010;
    16'b0100000000011000: out_v[390] = 10'b1011001100;
    16'b1100010010100000: out_v[390] = 10'b1101010100;
    default: out_v[390] = 10'd0;
  endcase
end

always @(*) begin
  case (addr)
    16'b0000010010000000: out_v[391] = 10'b0010110111;
    16'b0100010010010011: out_v[391] = 10'b1111001110;
    16'b0100011010010001: out_v[391] = 10'b0001111111;
    16'b0000011010000000: out_v[391] = 10'b1001110011;
    16'b0000011010010001: out_v[391] = 10'b0100010011;
    16'b0100110010010011: out_v[391] = 10'b0011101010;
    16'b0100000000010001: out_v[391] = 10'b1010111011;
    16'b0100001000010001: out_v[391] = 10'b0010011111;
    16'b0000000000010000: out_v[391] = 10'b0111110011;
    16'b0100110010010001: out_v[391] = 10'b0111101110;
    16'b0100011010010000: out_v[391] = 10'b1001111110;
    16'b0000010010010000: out_v[391] = 10'b1100110011;
    16'b0100010011010011: out_v[391] = 10'b1110111010;
    16'b0100010010010001: out_v[391] = 10'b0011101111;
    16'b1000011010010001: out_v[391] = 10'b1000010001;
    16'b0100011010010011: out_v[391] = 10'b0110110110;
    16'b1100011010010001: out_v[391] = 10'b1001010010;
    16'b0000011010010000: out_v[391] = 10'b1101110110;
    16'b1000001010010001: out_v[391] = 10'b0010011110;
    16'b1100001010010001: out_v[391] = 10'b0011101111;
    16'b0100010010010010: out_v[391] = 10'b1011001111;
    16'b0100111010010001: out_v[391] = 10'b1100111110;
    16'b0100001010010001: out_v[391] = 10'b1001101011;
    16'b1000011010000000: out_v[391] = 10'b0011000101;
    16'b0100010010000011: out_v[391] = 10'b0101011001;
    16'b1100001000010001: out_v[391] = 10'b1010010100;
    16'b0000010010010001: out_v[391] = 10'b1011000111;
    16'b0000010011010000: out_v[391] = 10'b0110111010;
    16'b0100001000000001: out_v[391] = 10'b1010011011;
    16'b0100011000010001: out_v[391] = 10'b1111001110;
    16'b0100010000010001: out_v[391] = 10'b1101111111;
    16'b0100011011010011: out_v[391] = 10'b1101010111;
    16'b1000011010010000: out_v[391] = 10'b0010110110;
    16'b0100010011010001: out_v[391] = 10'b1110110110;
    16'b0000011011010001: out_v[391] = 10'b0110110111;
    16'b0000000000000000: out_v[391] = 10'b0010011111;
    16'b0100010010010000: out_v[391] = 10'b1101101010;
    16'b0100010011000011: out_v[391] = 10'b1001111011;
    16'b0000010011010011: out_v[391] = 10'b1110101110;
    16'b0110010010010011: out_v[391] = 10'b1010111011;
    16'b0000010011010001: out_v[391] = 10'b0100110011;
    16'b0110010010010001: out_v[391] = 10'b1011100001;
    16'b0010000000011010: out_v[391] = 10'b0100100000;
    16'b0010000000001000: out_v[391] = 10'b1101010011;
    16'b0000000000001000: out_v[391] = 10'b1101001000;
    16'b0000000001001000: out_v[391] = 10'b1010101000;
    16'b0010000001001000: out_v[391] = 10'b1101100100;
    16'b0010000000000000: out_v[391] = 10'b1010010111;
    16'b0010000000001010: out_v[391] = 10'b0110101001;
    16'b0000000000011000: out_v[391] = 10'b0110110010;
    16'b0000000000011010: out_v[391] = 10'b1101000011;
    16'b0010000000011000: out_v[391] = 10'b1111111010;
    16'b0010000001011000: out_v[391] = 10'b0000110110;
    16'b0000000000001010: out_v[391] = 10'b1011001011;
    16'b1010000000011000: out_v[391] = 10'b1011101011;
    16'b0010001000000000: out_v[391] = 10'b0010010111;
    16'b1010001000011000: out_v[391] = 10'b1011101110;
    16'b0011000001011000: out_v[391] = 10'b1110001011;
    16'b1010001000001000: out_v[391] = 10'b0100001010;
    16'b1000000000011000: out_v[391] = 10'b0011100010;
    16'b0010001000001000: out_v[391] = 10'b1011011101;
    16'b0010000000011001: out_v[391] = 10'b1011010001;
    16'b0010001000011000: out_v[391] = 10'b1001110110;
    16'b0010010010011001: out_v[391] = 10'b1000011110;
    16'b0010010010011000: out_v[391] = 10'b1110000111;
    16'b0010001000011001: out_v[391] = 10'b0101011010;
    16'b1010001000000000: out_v[391] = 10'b1000100110;
    16'b0000001000001000: out_v[391] = 10'b1100100110;
    16'b0010000000001001: out_v[391] = 10'b0010111111;
    16'b0010011010010000: out_v[391] = 10'b1101010100;
    16'b0010001010011000: out_v[391] = 10'b1001101011;
    16'b1010001000010000: out_v[391] = 10'b0100101101;
    16'b0010000000010000: out_v[391] = 10'b1001111100;
    16'b0000001000011000: out_v[391] = 10'b0000110100;
    16'b1000001000011000: out_v[391] = 10'b1011110111;
    16'b1000000000001000: out_v[391] = 10'b1010001001;
    16'b1010000000001000: out_v[391] = 10'b0010100101;
    16'b0010001000010000: out_v[391] = 10'b0001001110;
    16'b1000001000001000: out_v[391] = 10'b0100100000;
    16'b0010011010011000: out_v[391] = 10'b1100000111;
    16'b0010011010011001: out_v[391] = 10'b1000101111;
    16'b0010010000011000: out_v[391] = 10'b1000110101;
    16'b1010001010011000: out_v[391] = 10'b1011111111;
    16'b0010000010011000: out_v[391] = 10'b0111101000;
    16'b0010010010010000: out_v[391] = 10'b0000101010;
    16'b0000011000000000: out_v[391] = 10'b0111011010;
    16'b1000000000000000: out_v[391] = 10'b0000110110;
    16'b0000011000011000: out_v[391] = 10'b0011011001;
    16'b0000011000001000: out_v[391] = 10'b0101101100;
    16'b0000001000010000: out_v[391] = 10'b1011111000;
    16'b0000010000000000: out_v[391] = 10'b0110001011;
    16'b0000001000000000: out_v[391] = 10'b0010100100;
    16'b1000011000010000: out_v[391] = 10'b1110001000;
    16'b0000011000010000: out_v[391] = 10'b1001001100;
    16'b1000011000001000: out_v[391] = 10'b0001110010;
    16'b1000010010010000: out_v[391] = 10'b1111011100;
    16'b0000010000010000: out_v[391] = 10'b1001101001;
    16'b0000000001000000: out_v[391] = 10'b1011000100;
    16'b0000011010001000: out_v[391] = 10'b1000101001;
    16'b1000010000000000: out_v[391] = 10'b0010111011;
    16'b0000010000001000: out_v[391] = 10'b0000111111;
    16'b1000010000010000: out_v[391] = 10'b0101111111;
    16'b1000011000000000: out_v[391] = 10'b0011100110;
    16'b1000011000011000: out_v[391] = 10'b0100110110;
    16'b0000010000011000: out_v[391] = 10'b1101001100;
    16'b0000011010011000: out_v[391] = 10'b1011010100;
    16'b0000000001010000: out_v[391] = 10'b1011101111;
    16'b0010001010001000: out_v[391] = 10'b0101111011;
    16'b0010011010001000: out_v[391] = 10'b1111110111;
    16'b0010001000001001: out_v[391] = 10'b0111001110;
    16'b0010000010001000: out_v[391] = 10'b1011111010;
    16'b0000010010001000: out_v[391] = 10'b1101010010;
    16'b0010010010001000: out_v[391] = 10'b1010101110;
    16'b0110010010001000: out_v[391] = 10'b1000110011;
    16'b0010010000001000: out_v[391] = 10'b0111110001;
    16'b0000000000001001: out_v[391] = 10'b1101100011;
    16'b0010000010001011: out_v[391] = 10'b1011011111;
    16'b0110011010001000: out_v[391] = 10'b1000011011;
    16'b0010011010001011: out_v[391] = 10'b1111111111;
    16'b0010010010001001: out_v[391] = 10'b0000101111;
    16'b0010010000001010: out_v[391] = 10'b1011111111;
    16'b0010000010001001: out_v[391] = 10'b1001011010;
    16'b0110010010001001: out_v[391] = 10'b1001010010;
    16'b0000010010001001: out_v[391] = 10'b1100100100;
    16'b0100010010001001: out_v[391] = 10'b1100011111;
    16'b0010011000001000: out_v[391] = 10'b0110000010;
    16'b0000011000001001: out_v[391] = 10'b1111001111;
    16'b0010010000001001: out_v[391] = 10'b0110110000;
    16'b0000011010001001: out_v[391] = 10'b1000111011;
    16'b0000000010001000: out_v[391] = 10'b0100110011;
    16'b0000001010001000: out_v[391] = 10'b0101011010;
    16'b0110011010001001: out_v[391] = 10'b1111010011;
    16'b0000010000001001: out_v[391] = 10'b0111011100;
    16'b0010000000000001: out_v[391] = 10'b0110011010;
    16'b0010000000001011: out_v[391] = 10'b1110101111;
    16'b0010000000000010: out_v[391] = 10'b0001111100;
    16'b0010010010001011: out_v[391] = 10'b1111101101;
    16'b0010011010001001: out_v[391] = 10'b1100111011;
    16'b0010010000001011: out_v[391] = 10'b1101100110;
    16'b0000011010001011: out_v[391] = 10'b0111111110;
    16'b0010011000001001: out_v[391] = 10'b1111011011;
    16'b0000001000001001: out_v[391] = 10'b1111100111;
    16'b0110000000011000: out_v[391] = 10'b0011110100;
    16'b0100000000011000: out_v[391] = 10'b1110110110;
    16'b0000000000000010: out_v[391] = 10'b1010110000;
    16'b0000000000010010: out_v[391] = 10'b0010110110;
    16'b0000001000001010: out_v[391] = 10'b0101010101;
    16'b0110000000001000: out_v[391] = 10'b1000100111;
    16'b0000001000010010: out_v[391] = 10'b1000010011;
    16'b0000001000000010: out_v[391] = 10'b0101100010;
    16'b0010001000001010: out_v[391] = 10'b1111010111;
    16'b1000001000000000: out_v[391] = 10'b1111000100;
    16'b0000001000011010: out_v[391] = 10'b1011111101;
    16'b0011010010001000: out_v[391] = 10'b1111000011;
    16'b0011000001000000: out_v[391] = 10'b1111001111;
    16'b0011010001001000: out_v[391] = 10'b0111101111;
    16'b0011000001001100: out_v[391] = 10'b1111011101;
    16'b0010010010000000: out_v[391] = 10'b1101101110;
    16'b0010010000000000: out_v[391] = 10'b0101010010;
    16'b0001010001001000: out_v[391] = 10'b1111100101;
    16'b0011000000000000: out_v[391] = 10'b0010111101;
    16'b0000000001001100: out_v[391] = 10'b0000101110;
    16'b0011000000001000: out_v[391] = 10'b1010001111;
    16'b0010000001001100: out_v[391] = 10'b1000110010;
    16'b0001000001001000: out_v[391] = 10'b0111010001;
    16'b0001010010001000: out_v[391] = 10'b1111101011;
    16'b0010011010000000: out_v[391] = 10'b1110100001;
    16'b0001000000001000: out_v[391] = 10'b1101000101;
    16'b0011010000001000: out_v[391] = 10'b0100001011;
    16'b0011010000000000: out_v[391] = 10'b0110100011;
    16'b0011000001001000: out_v[391] = 10'b0110100111;
    16'b0001000001001100: out_v[391] = 10'b0001010110;
    16'b0001010000001000: out_v[391] = 10'b1110011111;
    16'b0010011000000000: out_v[391] = 10'b1001011011;
    16'b0110011010000000: out_v[391] = 10'b0011111011;
    16'b0010000010000000: out_v[391] = 10'b1011000010;
    16'b0010001010000000: out_v[391] = 10'b0111001101;
    16'b0000001010000000: out_v[391] = 10'b0100011010;
    16'b0110000010000000: out_v[391] = 10'b0110011111;
    16'b0000011010000001: out_v[391] = 10'b0111001110;
    16'b0100011010000000: out_v[391] = 10'b0111000110;
    16'b0110010010000000: out_v[391] = 10'b0011011000;
    16'b0000000010000000: out_v[391] = 10'b0110100010;
    16'b0110001010000000: out_v[391] = 10'b0111110010;
    16'b0100011010000001: out_v[391] = 10'b0111001110;
    16'b0100010010000000: out_v[391] = 10'b1011001011;
    16'b0000011010100000: out_v[391] = 10'b1111111111;
    16'b0110001010001000: out_v[391] = 10'b0100011110;
    16'b0100000010011000: out_v[391] = 10'b0101011001;
    16'b0110010010011000: out_v[391] = 10'b0110000110;
    16'b0110000010011010: out_v[391] = 10'b0110101100;
    16'b0110001010011000: out_v[391] = 10'b1101100001;
    16'b0110000010011000: out_v[391] = 10'b0010111110;
    16'b0010000001011010: out_v[391] = 10'b1110111010;
    16'b0010000010011010: out_v[391] = 10'b0100011111;
    16'b0110001010011010: out_v[391] = 10'b0111101011;
    16'b0100001010011000: out_v[391] = 10'b0110010010;
    16'b0110011010011000: out_v[391] = 10'b0111100110;
    16'b0110000010001000: out_v[391] = 10'b0111000101;
    16'b0010001000011010: out_v[391] = 10'b1100110001;
    16'b0000001010011000: out_v[391] = 10'b0101110011;
    16'b0010011010000001: out_v[391] = 10'b1001100010;
    16'b1010011010001001: out_v[391] = 10'b0011101111;
    16'b1000011010001001: out_v[391] = 10'b1101100111;
    16'b0000000010001001: out_v[391] = 10'b1101100011;
    default: out_v[391] = 10'd0;
  endcase
end


endmodule